library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.ALL;

entity ROM_1 is
    Port ( addr : in STD_LOGIC_VECTOR (11 downto 0);
           Cout : out STD_LOGIC_VECTOR (19 downto 0));
end ROM_1;

architecture Behavioral of ROM_1 is
type vector is Array(0 to 4095) of Std_logic_vector(19 downto 0);
Constant memory: vector:=
(0=>x"00064",
1=>x"00063",
2=>x"00062",
3=>x"00061",
4=>x"00060",
5=>x"0005f",
6=>x"0005e",
7=>x"0005d",
8=>x"0005c",
9=>x"0005b",
10=>x"0005a",
11=>x"0005a",
12=>x"00059",
13=>x"00058",
14=>x"00057",
15=>x"00056",
16=>x"00056",
17=>x"00055",
18=>x"00054",
19=>x"00054",
20=>x"00053",
21=>x"00052",
22=>x"00051",
23=>x"00051",
24=>x"00050",
25=>x"00050",
26=>x"0004f",
27=>x"0004e",
28=>x"0004e",
29=>x"0004d",
30=>x"0004c",
31=>x"0004c",
32=>x"0004b",
33=>x"0004b",
34=>x"0004a",
35=>x"0004a",
36=>x"00049",
37=>x"00048",
38=>x"00048",
39=>x"00047",
40=>x"00047",
41=>x"00046",
42=>x"00046",
43=>x"00045",
44=>x"00045",
45=>x"00044",
46=>x"00044",
47=>x"00044",
48=>x"00043",
49=>x"00043",
50=>x"00042",
51=>x"00042",
52=>x"00041",
53=>x"00041",
54=>x"00040",
55=>x"00040",
56=>x"00040",
57=>x"0003f",
58=>x"0003f",
59=>x"0003e",
60=>x"0003e",
61=>x"0003e",
62=>x"0003d",
63=>x"0003d",
64=>x"0003c",
65=>x"0003c",
66=>x"0003c",
67=>x"0003b",
68=>x"0003b",
69=>x"0003b",
70=>x"0003a",
71=>x"0003a",
72=>x"0003a",
73=>x"00039",
74=>x"00039",
75=>x"00039",
76=>x"00038",
77=>x"00038",
78=>x"00038",
79=>x"00037",
80=>x"00037",
81=>x"00037",
82=>x"00036",
83=>x"00036",
84=>x"00036",
85=>x"00036",
86=>x"00035",
87=>x"00035",
88=>x"00035",
89=>x"00034",
90=>x"00034",
91=>x"00034",
92=>x"00034",
93=>x"00033",
94=>x"00033",
95=>x"00033",
96=>x"00033",
97=>x"00032",
98=>x"00032",
99=>x"00032",
100=>x"00032",
101=>x"00031",
102=>x"00031",
103=>x"00031",
104=>x"00031",
105=>x"00030",
106=>x"00030",
107=>x"00030",
108=>x"00030",
109=>x"0002f",
110=>x"0002f",
111=>x"0002f",
112=>x"0002f",
113=>x"0002e",
114=>x"0002e",
115=>x"0002e",
116=>x"0002e",
117=>x"0002e",
118=>x"0002d",
119=>x"0002d",
120=>x"0002d",
121=>x"0002d",
122=>x"0002d",
123=>x"0002c",
124=>x"0002c",
125=>x"0002c",
126=>x"0002c",
127=>x"0002c",
128=>x"0002b",
129=>x"0002b",
130=>x"0002b",
131=>x"0002b",
132=>x"0002b",
133=>x"0002a",
134=>x"0002a",
135=>x"0002a",
136=>x"0002a",
137=>x"0002a",
138=>x"0002a",
139=>x"00029",
140=>x"00029",
141=>x"00029",
142=>x"00029",
143=>x"00029",
144=>x"00028",
145=>x"00028",
146=>x"00028",
147=>x"00028",
148=>x"00028",
149=>x"00028",
150=>x"00028",
151=>x"00027",
152=>x"00027",
153=>x"00027",
154=>x"00027",
155=>x"00027",
156=>x"00027",
157=>x"00026",
158=>x"00026",
159=>x"00026",
160=>x"00026",
161=>x"00026",
162=>x"00026",
163=>x"00026",
164=>x"00025",
165=>x"00025",
166=>x"00025",
167=>x"00025",
168=>x"00025",
169=>x"00025",
170=>x"00025",
171=>x"00024",
172=>x"00024",
173=>x"00024",
174=>x"00024",
175=>x"00024",
176=>x"00024",
177=>x"00024",
178=>x"00023",
179=>x"00023",
180=>x"00023",
181=>x"00023",
182=>x"00023",
183=>x"00023",
184=>x"00023",
185=>x"00023",
186=>x"00022",
187=>x"00022",
188=>x"00022",
189=>x"00022",
190=>x"00022",
191=>x"00022",
192=>x"00022",
193=>x"00022",
194=>x"00022",
195=>x"00021",
196=>x"00021",
197=>x"00021",
198=>x"00021",
199=>x"00021",
200=>x"00021",
201=>x"00021",
202=>x"00021",
203=>x"00021",
204=>x"00020",
205=>x"00020",
206=>x"00020",
207=>x"00020",
208=>x"00020",
209=>x"00020",
210=>x"00020",
211=>x"00020",
212=>x"00020",
213=>x"0001f",
214=>x"0001f",
215=>x"0001f",
216=>x"0001f",
217=>x"0001f",
218=>x"0001f",
219=>x"0001f",
220=>x"0001f",
221=>x"0001f",
222=>x"0001f",
223=>x"0001e",
224=>x"0001e",
225=>x"0001e",
226=>x"0001e",
227=>x"0001e",
228=>x"0001e",
229=>x"0001e",
230=>x"0001e",
231=>x"0001e",
232=>x"0001e",
233=>x"0001e",
234=>x"0001d",
235=>x"0001d",
236=>x"0001d",
237=>x"0001d",
238=>x"0001d",
239=>x"0001d",
240=>x"0001d",
241=>x"0001d",
242=>x"0001d",
243=>x"0001d",
244=>x"0001d",
245=>x"0001c",
246=>x"0001c",
247=>x"0001c",
248=>x"0001c",
249=>x"0001c",
250=>x"0001c",
251=>x"0001c",
252=>x"0001c",
253=>x"0001c",
254=>x"0001c",
255=>x"0001c",
256=>x"0001c",
257=>x"0001c",
258=>x"0001b",
259=>x"0001b",
260=>x"0001b",
261=>x"0001b",
262=>x"0001b",
263=>x"0001b",
264=>x"0001b",
265=>x"0001b",
266=>x"0001b",
267=>x"0001b",
268=>x"0001b",
269=>x"0001b",
270=>x"0001b",
271=>x"0001a",
272=>x"0001a",
273=>x"0001a",
274=>x"0001a",
275=>x"0001a",
276=>x"0001a",
277=>x"0001a",
278=>x"0001a",
279=>x"0001a",
280=>x"0001a",
281=>x"0001a",
282=>x"0001a",
283=>x"0001a",
284=>x"0001a",
285=>x"00019",
286=>x"00019",
287=>x"00019",
288=>x"00019",
289=>x"00019",
290=>x"00019",
291=>x"00019",
292=>x"00019",
293=>x"00019",
294=>x"00019",
295=>x"00019",
296=>x"00019",
297=>x"00019",
298=>x"00019",
299=>x"00019",
300=>x"00019",
301=>x"00018",
302=>x"00018",
303=>x"00018",
304=>x"00018",
305=>x"00018",
306=>x"00018",
307=>x"00018",
308=>x"00018",
309=>x"00018",
310=>x"00018",
311=>x"00018",
312=>x"00018",
313=>x"00018",
314=>x"00018",
315=>x"00018",
316=>x"00018",
317=>x"00017",
318=>x"00017",
319=>x"00017",
320=>x"00017",
321=>x"00017",
322=>x"00017",
323=>x"00017",
324=>x"00017",
325=>x"00017",
326=>x"00017",
327=>x"00017",
328=>x"00017",
329=>x"00017",
330=>x"00017",
331=>x"00017",
332=>x"00017",
333=>x"00017",
334=>x"00017",
335=>x"00016",
336=>x"00016",
337=>x"00016",
338=>x"00016",
339=>x"00016",
340=>x"00016",
341=>x"00016",
342=>x"00016",
343=>x"00016",
344=>x"00016",
345=>x"00016",
346=>x"00016",
347=>x"00016",
348=>x"00016",
349=>x"00016",
350=>x"00016",
351=>x"00016",
352=>x"00016",
353=>x"00016",
354=>x"00016",
355=>x"00015",
356=>x"00015",
357=>x"00015",
358=>x"00015",
359=>x"00015",
360=>x"00015",
361=>x"00015",
362=>x"00015",
363=>x"00015",
364=>x"00015",
365=>x"00015",
366=>x"00015",
367=>x"00015",
368=>x"00015",
369=>x"00015",
370=>x"00015",
371=>x"00015",
372=>x"00015",
373=>x"00015",
374=>x"00015",
375=>x"00015",
376=>x"00015",
377=>x"00014",
378=>x"00014",
379=>x"00014",
380=>x"00014",
381=>x"00014",
382=>x"00014",
383=>x"00014",
384=>x"00014",
385=>x"00014",
386=>x"00014",
387=>x"00014",
388=>x"00014",
389=>x"00014",
390=>x"00014",
391=>x"00014",
392=>x"00014",
393=>x"00014",
394=>x"00014",
395=>x"00014",
396=>x"00014",
397=>x"00014",
398=>x"00014",
399=>x"00014",
400=>x"00014",
401=>x"00013",
402=>x"00013",
403=>x"00013",
404=>x"00013",
405=>x"00013",
406=>x"00013",
407=>x"00013",
408=>x"00013",
409=>x"00013",
410=>x"00013",
411=>x"00013",
412=>x"00013",
413=>x"00013",
414=>x"00013",
415=>x"00013",
416=>x"00013",
417=>x"00013",
418=>x"00013",
419=>x"00013",
420=>x"00013",
421=>x"00013",
422=>x"00013",
423=>x"00013",
424=>x"00013",
425=>x"00013",
426=>x"00013",
427=>x"00012",
428=>x"00012",
429=>x"00012",
430=>x"00012",
431=>x"00012",
432=>x"00012",
433=>x"00012",
434=>x"00012",
435=>x"00012",
436=>x"00012",
437=>x"00012",
438=>x"00012",
439=>x"00012",
440=>x"00012",
441=>x"00012",
442=>x"00012",
443=>x"00012",
444=>x"00012",
445=>x"00012",
446=>x"00012",
447=>x"00012",
448=>x"00012",
449=>x"00012",
450=>x"00012",
451=>x"00012",
452=>x"00012",
453=>x"00012",
454=>x"00012",
455=>x"00012",
456=>x"00011",
457=>x"00011",
458=>x"00011",
459=>x"00011",
460=>x"00011",
461=>x"00011",
462=>x"00011",
463=>x"00011",
464=>x"00011",
465=>x"00011",
466=>x"00011",
467=>x"00011",
468=>x"00011",
469=>x"00011",
470=>x"00011",
471=>x"00011",
472=>x"00011",
473=>x"00011",
474=>x"00011",
475=>x"00011",
476=>x"00011",
477=>x"00011",
478=>x"00011",
479=>x"00011",
480=>x"00011",
481=>x"00011",
482=>x"00011",
483=>x"00011",
484=>x"00011",
485=>x"00011",
486=>x"00011",
487=>x"00011",
488=>x"00011",
489=>x"00010",
490=>x"00010",
491=>x"00010",
492=>x"00010",
493=>x"00010",
494=>x"00010",
495=>x"00010",
496=>x"00010",
497=>x"00010",
498=>x"00010",
499=>x"00010",
500=>x"00010",
501=>x"00010",
502=>x"00010",
503=>x"00010",
504=>x"00010",
505=>x"00010",
506=>x"00010",
507=>x"00010",
508=>x"00010",
509=>x"00010",
510=>x"00010",
511=>x"00010",
512=>x"00010",
513=>x"00010",
514=>x"00010",
515=>x"00010",
516=>x"00010",
517=>x"00010",
518=>x"00010",
519=>x"00010",
520=>x"00010",
521=>x"00010",
522=>x"00010",
523=>x"00010",
524=>x"00010",
525=>x"00010",
526=>x"0000f",
527=>x"0000f",
528=>x"0000f",
529=>x"0000f",
530=>x"0000f",
531=>x"0000f",
532=>x"0000f",
533=>x"0000f",
534=>x"0000f",
535=>x"0000f",
536=>x"0000f",
537=>x"0000f",
538=>x"0000f",
539=>x"0000f",
540=>x"0000f",
541=>x"0000f",
542=>x"0000f",
543=>x"0000f",
544=>x"0000f",
545=>x"0000f",
546=>x"0000f",
547=>x"0000f",
548=>x"0000f",
549=>x"0000f",
550=>x"0000f",
551=>x"0000f",
552=>x"0000f",
553=>x"0000f",
554=>x"0000f",
555=>x"0000f",
556=>x"0000f",
557=>x"0000f",
558=>x"0000f",
559=>x"0000f",
560=>x"0000f",
561=>x"0000f",
562=>x"0000f",
563=>x"0000f",
564=>x"0000f",
565=>x"0000f",
566=>x"0000f",
567=>x"0000e",
568=>x"0000e",
569=>x"0000e",
570=>x"0000e",
571=>x"0000e",
572=>x"0000e",
573=>x"0000e",
574=>x"0000e",
575=>x"0000e",
576=>x"0000e",
577=>x"0000e",
578=>x"0000e",
579=>x"0000e",
580=>x"0000e",
581=>x"0000e",
582=>x"0000e",
583=>x"0000e",
584=>x"0000e",
585=>x"0000e",
586=>x"0000e",
587=>x"0000e",
588=>x"0000e",
589=>x"0000e",
590=>x"0000e",
591=>x"0000e",
592=>x"0000e",
593=>x"0000e",
594=>x"0000e",
595=>x"0000e",
596=>x"0000e",
597=>x"0000e",
598=>x"0000e",
599=>x"0000e",
600=>x"0000e",
601=>x"0000e",
602=>x"0000e",
603=>x"0000e",
604=>x"0000e",
605=>x"0000e",
606=>x"0000e",
607=>x"0000e",
608=>x"0000e",
609=>x"0000e",
610=>x"0000e",
611=>x"0000e",
612=>x"0000e",
613=>x"0000e",
614=>x"0000e",
615=>x"0000d",
616=>x"0000d",
617=>x"0000d",
618=>x"0000d",
619=>x"0000d",
620=>x"0000d",
621=>x"0000d",
622=>x"0000d",
623=>x"0000d",
624=>x"0000d",
625=>x"0000d",
626=>x"0000d",
627=>x"0000d",
628=>x"0000d",
629=>x"0000d",
630=>x"0000d",
631=>x"0000d",
632=>x"0000d",
633=>x"0000d",
634=>x"0000d",
635=>x"0000d",
636=>x"0000d",
637=>x"0000d",
638=>x"0000d",
639=>x"0000d",
640=>x"0000d",
641=>x"0000d",
642=>x"0000d",
643=>x"0000d",
644=>x"0000d",
645=>x"0000d",
646=>x"0000d",
647=>x"0000d",
648=>x"0000d",
649=>x"0000d",
650=>x"0000d",
651=>x"0000d",
652=>x"0000d",
653=>x"0000d",
654=>x"0000d",
655=>x"0000d",
656=>x"0000d",
657=>x"0000d",
658=>x"0000d",
659=>x"0000d",
660=>x"0000d",
661=>x"0000d",
662=>x"0000d",
663=>x"0000d",
664=>x"0000d",
665=>x"0000d",
666=>x"0000d",
667=>x"0000d",
668=>x"0000d",
669=>x"0000d",
670=>x"0000c",
671=>x"0000c",
672=>x"0000c",
673=>x"0000c",
674=>x"0000c",
675=>x"0000c",
676=>x"0000c",
677=>x"0000c",
678=>x"0000c",
679=>x"0000c",
680=>x"0000c",
681=>x"0000c",
682=>x"0000c",
683=>x"0000c",
684=>x"0000c",
685=>x"0000c",
686=>x"0000c",
687=>x"0000c",
688=>x"0000c",
689=>x"0000c",
690=>x"0000c",
691=>x"0000c",
692=>x"0000c",
693=>x"0000c",
694=>x"0000c",
695=>x"0000c",
696=>x"0000c",
697=>x"0000c",
698=>x"0000c",
699=>x"0000c",
700=>x"0000c",
701=>x"0000c",
702=>x"0000c",
703=>x"0000c",
704=>x"0000c",
705=>x"0000c",
706=>x"0000c",
707=>x"0000c",
708=>x"0000c",
709=>x"0000c",
710=>x"0000c",
711=>x"0000c",
712=>x"0000c",
713=>x"0000c",
714=>x"0000c",
715=>x"0000c",
716=>x"0000c",
717=>x"0000c",
718=>x"0000c",
719=>x"0000c",
720=>x"0000c",
721=>x"0000c",
722=>x"0000c",
723=>x"0000c",
724=>x"0000c",
725=>x"0000c",
726=>x"0000c",
727=>x"0000c",
728=>x"0000c",
729=>x"0000c",
730=>x"0000c",
731=>x"0000c",
732=>x"0000c",
733=>x"0000c",
734=>x"0000b",
735=>x"0000b",
736=>x"0000b",
737=>x"0000b",
738=>x"0000b",
739=>x"0000b",
740=>x"0000b",
741=>x"0000b",
742=>x"0000b",
743=>x"0000b",
744=>x"0000b",
745=>x"0000b",
746=>x"0000b",
747=>x"0000b",
748=>x"0000b",
749=>x"0000b",
750=>x"0000b",
751=>x"0000b",
752=>x"0000b",
753=>x"0000b",
754=>x"0000b",
755=>x"0000b",
756=>x"0000b",
757=>x"0000b",
758=>x"0000b",
759=>x"0000b",
760=>x"0000b",
761=>x"0000b",
762=>x"0000b",
763=>x"0000b",
764=>x"0000b",
765=>x"0000b",
766=>x"0000b",
767=>x"0000b",
768=>x"0000b",
769=>x"0000b",
770=>x"0000b",
771=>x"0000b",
772=>x"0000b",
773=>x"0000b",
774=>x"0000b",
775=>x"0000b",
776=>x"0000b",
777=>x"0000b",
778=>x"0000b",
779=>x"0000b",
780=>x"0000b",
781=>x"0000b",
782=>x"0000b",
783=>x"0000b",
784=>x"0000b",
785=>x"0000b",
786=>x"0000b",
787=>x"0000b",
788=>x"0000b",
789=>x"0000b",
790=>x"0000b",
791=>x"0000b",
792=>x"0000b",
793=>x"0000b",
794=>x"0000b",
795=>x"0000b",
796=>x"0000b",
797=>x"0000b",
798=>x"0000b",
799=>x"0000b",
800=>x"0000b",
801=>x"0000b",
802=>x"0000b",
803=>x"0000b",
804=>x"0000b",
805=>x"0000b",
806=>x"0000b",
807=>x"0000b",
808=>x"0000b",
809=>x"0000b",
810=>x"0000a",
811=>x"0000a",
812=>x"0000a",
813=>x"0000a",
814=>x"0000a",
815=>x"0000a",
816=>x"0000a",
817=>x"0000a",
818=>x"0000a",
819=>x"0000a",
820=>x"0000a",
821=>x"0000a",
822=>x"0000a",
823=>x"0000a",
824=>x"0000a",
825=>x"0000a",
826=>x"0000a",
827=>x"0000a",
828=>x"0000a",
829=>x"0000a",
830=>x"0000a",
831=>x"0000a",
832=>x"0000a",
833=>x"0000a",
834=>x"0000a",
835=>x"0000a",
836=>x"0000a",
837=>x"0000a",
838=>x"0000a",
839=>x"0000a",
840=>x"0000a",
841=>x"0000a",
842=>x"0000a",
843=>x"0000a",
844=>x"0000a",
845=>x"0000a",
846=>x"0000a",
847=>x"0000a",
848=>x"0000a",
849=>x"0000a",
850=>x"0000a",
851=>x"0000a",
852=>x"0000a",
853=>x"0000a",
854=>x"0000a",
855=>x"0000a",
856=>x"0000a",
857=>x"0000a",
858=>x"0000a",
859=>x"0000a",
860=>x"0000a",
861=>x"0000a",
862=>x"0000a",
863=>x"0000a",
864=>x"0000a",
865=>x"0000a",
866=>x"0000a",
867=>x"0000a",
868=>x"0000a",
869=>x"0000a",
870=>x"0000a",
871=>x"0000a",
872=>x"0000a",
873=>x"0000a",
874=>x"0000a",
875=>x"0000a",
876=>x"0000a",
877=>x"0000a",
878=>x"0000a",
879=>x"0000a",
880=>x"0000a",
881=>x"0000a",
882=>x"0000a",
883=>x"0000a",
884=>x"0000a",
885=>x"0000a",
886=>x"0000a",
887=>x"0000a",
888=>x"0000a",
889=>x"0000a",
890=>x"0000a",
891=>x"0000a",
892=>x"0000a",
893=>x"0000a",
894=>x"0000a",
895=>x"0000a",
896=>x"0000a",
897=>x"0000a",
898=>x"0000a",
899=>x"0000a",
900=>x"0000a",
901=>x"00009",
902=>x"00009",
903=>x"00009",
904=>x"00009",
905=>x"00009",
906=>x"00009",
907=>x"00009",
908=>x"00009",
909=>x"00009",
910=>x"00009",
911=>x"00009",
912=>x"00009",
913=>x"00009",
914=>x"00009",
915=>x"00009",
916=>x"00009",
917=>x"00009",
918=>x"00009",
919=>x"00009",
920=>x"00009",
921=>x"00009",
922=>x"00009",
923=>x"00009",
924=>x"00009",
925=>x"00009",
926=>x"00009",
927=>x"00009",
928=>x"00009",
929=>x"00009",
930=>x"00009",
931=>x"00009",
932=>x"00009",
933=>x"00009",
934=>x"00009",
935=>x"00009",
936=>x"00009",
937=>x"00009",
938=>x"00009",
939=>x"00009",
940=>x"00009",
941=>x"00009",
942=>x"00009",
943=>x"00009",
944=>x"00009",
945=>x"00009",
946=>x"00009",
947=>x"00009",
948=>x"00009",
949=>x"00009",
950=>x"00009",
951=>x"00009",
952=>x"00009",
953=>x"00009",
954=>x"00009",
955=>x"00009",
956=>x"00009",
957=>x"00009",
958=>x"00009",
959=>x"00009",
960=>x"00009",
961=>x"00009",
962=>x"00009",
963=>x"00009",
964=>x"00009",
965=>x"00009",
966=>x"00009",
967=>x"00009",
968=>x"00009",
969=>x"00009",
970=>x"00009",
971=>x"00009",
972=>x"00009",
973=>x"00009",
974=>x"00009",
975=>x"00009",
976=>x"00009",
977=>x"00009",
978=>x"00009",
979=>x"00009",
980=>x"00009",
981=>x"00009",
982=>x"00009",
983=>x"00009",
984=>x"00009",
985=>x"00009",
986=>x"00009",
987=>x"00009",
988=>x"00009",
989=>x"00009",
990=>x"00009",
991=>x"00009",
992=>x"00009",
993=>x"00009",
994=>x"00009",
995=>x"00009",
996=>x"00009",
997=>x"00009",
998=>x"00009",
999=>x"00009",
others=>x"00000"
);
begin
Cout<=memory(to_integer(unsigned(addr)));

end Behavioral;