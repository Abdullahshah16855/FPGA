library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.ALL;

entity ROM_128 is
    Port ( addr : in STD_LOGIC_VECTOR (11 downto 0);
           Cout : out STD_LOGIC_VECTOR (19 downto 0));
end ROM_128;

architecture Behavioral of ROM_128 is
type vector is Array(0 to 4095) of Std_logic_vector(19 downto 0);
Constant memory: vector:=
(
0=>x"00064",
1=>x"00063",
2=>x"00062",
3=>x"00061",
4=>x"00060",
5=>x"00060",
6=>x"0005f",
7=>x"0005e",
8=>x"0005e",
9=>x"0005d",
10=>x"0005c",
11=>x"0005c",
12=>x"0005b",
13=>x"0005a",
14=>x"0005a",
15=>x"00059",
16=>x"00058",
17=>x"00058",
18=>x"00057",
19=>x"00057",
20=>x"00056",
21=>x"00055",
22=>x"00055",
23=>x"00054",
24=>x"00054",
25=>x"00053",
26=>x"00053",
27=>x"00052",
28=>x"00052",
29=>x"00051",
30=>x"00051",
31=>x"00050",
32=>x"00050",
33=>x"0004f",
34=>x"0004f",
35=>x"0004e",
36=>x"0004e",
37=>x"0004d",
38=>x"0004d",
39=>x"0004c",
40=>x"0004c",
41=>x"0004b",
42=>x"0004b",
43=>x"0004a",
44=>x"0004a",
45=>x"00049",
46=>x"00049",
47=>x"00049",
48=>x"00048",
49=>x"00048",
50=>x"00047",
51=>x"00047",
52=>x"00047",
53=>x"00046",
54=>x"00046",
55=>x"00045",
56=>x"00045",
57=>x"00045",
58=>x"00044",
59=>x"00044",
60=>x"00044",
61=>x"00043",
62=>x"00043",
63=>x"00043",
64=>x"00042",
65=>x"00042",
66=>x"00041",
67=>x"00041",
68=>x"00041",
69=>x"00040",
70=>x"00040",
71=>x"00040",
72=>x"00040",
73=>x"0003f",
74=>x"0003f",
75=>x"0003f",
76=>x"0003e",
77=>x"0003e",
78=>x"0003e",
79=>x"0003d",
80=>x"0003d",
81=>x"0003d",
82=>x"0003c",
83=>x"0003c",
84=>x"0003c",
85=>x"0003c",
86=>x"0003b",
87=>x"0003b",
88=>x"0003b",
89=>x"0003a",
90=>x"0003a",
91=>x"0003a",
92=>x"0003a",
93=>x"00039",
94=>x"00039",
95=>x"00039",
96=>x"00039",
97=>x"00038",
98=>x"00038",
99=>x"00038",
100=>x"00038",
101=>x"00037",
102=>x"00037",
103=>x"00037",
104=>x"00037",
105=>x"00036",
106=>x"00036",
107=>x"00036",
108=>x"00036",
109=>x"00036",
110=>x"00035",
111=>x"00035",
112=>x"00035",
113=>x"00035",
114=>x"00034",
115=>x"00034",
116=>x"00034",
117=>x"00034",
118=>x"00034",
119=>x"00033",
120=>x"00033",
121=>x"00033",
122=>x"00033",
123=>x"00032",
124=>x"00032",
125=>x"00032",
126=>x"00032",
127=>x"00032",
128=>x"00032",
129=>x"00031",
130=>x"00031",
131=>x"00031",
132=>x"00031",
133=>x"00031",
134=>x"00030",
135=>x"00030",
136=>x"00030",
137=>x"00030",
138=>x"00030",
139=>x"0002f",
140=>x"0002f",
141=>x"0002f",
142=>x"0002f",
143=>x"0002f",
144=>x"0002f",
145=>x"0002e",
146=>x"0002e",
147=>x"0002e",
148=>x"0002e",
149=>x"0002e",
150=>x"0002e",
151=>x"0002d",
152=>x"0002d",
153=>x"0002d",
154=>x"0002d",
155=>x"0002d",
156=>x"0002d",
157=>x"0002c",
158=>x"0002c",
159=>x"0002c",
160=>x"0002c",
161=>x"0002c",
162=>x"0002c",
163=>x"0002b",
164=>x"0002b",
165=>x"0002b",
166=>x"0002b",
167=>x"0002b",
168=>x"0002b",
169=>x"0002b",
170=>x"0002a",
171=>x"0002a",
172=>x"0002a",
173=>x"0002a",
174=>x"0002a",
175=>x"0002a",
176=>x"0002a",
177=>x"00029",
178=>x"00029",
179=>x"00029",
180=>x"00029",
181=>x"00029",
182=>x"00029",
183=>x"00029",
184=>x"00029",
185=>x"00028",
186=>x"00028",
187=>x"00028",
188=>x"00028",
189=>x"00028",
190=>x"00028",
191=>x"00028",
192=>x"00028",
193=>x"00027",
194=>x"00027",
195=>x"00027",
196=>x"00027",
197=>x"00027",
198=>x"00027",
199=>x"00027",
200=>x"00027",
201=>x"00026",
202=>x"00026",
203=>x"00026",
204=>x"00026",
205=>x"00026",
206=>x"00026",
207=>x"00026",
208=>x"00026",
209=>x"00025",
210=>x"00025",
211=>x"00025",
212=>x"00025",
213=>x"00025",
214=>x"00025",
215=>x"00025",
216=>x"00025",
217=>x"00025",
218=>x"00024",
219=>x"00024",
220=>x"00024",
221=>x"00024",
222=>x"00024",
223=>x"00024",
224=>x"00024",
225=>x"00024",
226=>x"00024",
227=>x"00024",
228=>x"00023",
229=>x"00023",
230=>x"00023",
231=>x"00023",
232=>x"00023",
233=>x"00023",
234=>x"00023",
235=>x"00023",
236=>x"00023",
237=>x"00023",
238=>x"00022",
239=>x"00022",
240=>x"00022",
241=>x"00022",
242=>x"00022",
243=>x"00022",
244=>x"00022",
245=>x"00022",
246=>x"00022",
247=>x"00022",
248=>x"00022",
249=>x"00021",
250=>x"00021",
251=>x"00021",
252=>x"00021",
253=>x"00021",
254=>x"00021",
255=>x"00021",
256=>x"00021",
257=>x"00021",
258=>x"00021",
259=>x"00021",
260=>x"00020",
261=>x"00020",
262=>x"00020",
263=>x"00020",
264=>x"00020",
265=>x"00020",
266=>x"00020",
267=>x"00020",
268=>x"00020",
269=>x"00020",
270=>x"00020",
271=>x"00020",
272=>x"00020",
273=>x"0001f",
274=>x"0001f",
275=>x"0001f",
276=>x"0001f",
277=>x"0001f",
278=>x"0001f",
279=>x"0001f",
280=>x"0001f",
281=>x"0001f",
282=>x"0001f",
283=>x"0001f",
284=>x"0001f",
285=>x"0001e",
286=>x"0001e",
287=>x"0001e",
288=>x"0001e",
289=>x"0001e",
290=>x"0001e",
291=>x"0001e",
292=>x"0001e",
293=>x"0001e",
294=>x"0001e",
295=>x"0001e",
296=>x"0001e",
297=>x"0001e",
298=>x"0001e",
299=>x"0001d",
300=>x"0001d",
301=>x"0001d",
302=>x"0001d",
303=>x"0001d",
304=>x"0001d",
305=>x"0001d",
306=>x"0001d",
307=>x"0001d",
308=>x"0001d",
309=>x"0001d",
310=>x"0001d",
311=>x"0001d",
312=>x"0001d",
313=>x"0001d",
314=>x"0001c",
315=>x"0001c",
316=>x"0001c",
317=>x"0001c",
318=>x"0001c",
319=>x"0001c",
320=>x"0001c",
321=>x"0001c",
322=>x"0001c",
323=>x"0001c",
324=>x"0001c",
325=>x"0001c",
326=>x"0001c",
327=>x"0001c",
328=>x"0001c",
329=>x"0001c",
330=>x"0001b",
331=>x"0001b",
332=>x"0001b",
333=>x"0001b",
334=>x"0001b",
335=>x"0001b",
336=>x"0001b",
337=>x"0001b",
338=>x"0001b",
339=>x"0001b",
340=>x"0001b",
341=>x"0001b",
342=>x"0001b",
343=>x"0001b",
344=>x"0001b",
345=>x"0001b",
346=>x"0001b",
347=>x"0001a",
348=>x"0001a",
349=>x"0001a",
350=>x"0001a",
351=>x"0001a",
352=>x"0001a",
353=>x"0001a",
354=>x"0001a",
355=>x"0001a",
356=>x"0001a",
357=>x"0001a",
358=>x"0001a",
359=>x"0001a",
360=>x"0001a",
361=>x"0001a",
362=>x"0001a",
363=>x"0001a",
364=>x"0001a",
365=>x"00019",
366=>x"00019",
367=>x"00019",
368=>x"00019",
369=>x"00019",
370=>x"00019",
371=>x"00019",
372=>x"00019",
373=>x"00019",
374=>x"00019",
375=>x"00019",
376=>x"00019",
377=>x"00019",
378=>x"00019",
379=>x"00019",
380=>x"00019",
381=>x"00019",
382=>x"00019",
383=>x"00019",
384=>x"00019",
385=>x"00018",
386=>x"00018",
387=>x"00018",
388=>x"00018",
389=>x"00018",
390=>x"00018",
391=>x"00018",
392=>x"00018",
393=>x"00018",
394=>x"00018",
395=>x"00018",
396=>x"00018",
397=>x"00018",
398=>x"00018",
399=>x"00018",
400=>x"00018",
401=>x"00018",
402=>x"00018",
403=>x"00018",
404=>x"00018",
405=>x"00018",
406=>x"00017",
407=>x"00017",
408=>x"00017",
409=>x"00017",
410=>x"00017",
411=>x"00017",
412=>x"00017",
413=>x"00017",
414=>x"00017",
415=>x"00017",
416=>x"00017",
417=>x"00017",
418=>x"00017",
419=>x"00017",
420=>x"00017",
421=>x"00017",
422=>x"00017",
423=>x"00017",
424=>x"00017",
425=>x"00017",
426=>x"00017",
427=>x"00017",
428=>x"00017",
429=>x"00016",
430=>x"00016",
431=>x"00016",
432=>x"00016",
433=>x"00016",
434=>x"00016",
435=>x"00016",
436=>x"00016",
437=>x"00016",
438=>x"00016",
439=>x"00016",
440=>x"00016",
441=>x"00016",
442=>x"00016",
443=>x"00016",
444=>x"00016",
445=>x"00016",
446=>x"00016",
447=>x"00016",
448=>x"00016",
449=>x"00016",
450=>x"00016",
451=>x"00016",
452=>x"00016",
453=>x"00016",
454=>x"00015",
455=>x"00015",
456=>x"00015",
457=>x"00015",
458=>x"00015",
459=>x"00015",
460=>x"00015",
461=>x"00015",
462=>x"00015",
463=>x"00015",
464=>x"00015",
465=>x"00015",
466=>x"00015",
467=>x"00015",
468=>x"00015",
469=>x"00015",
470=>x"00015",
471=>x"00015",
472=>x"00015",
473=>x"00015",
474=>x"00015",
475=>x"00015",
476=>x"00015",
477=>x"00015",
478=>x"00015",
479=>x"00015",
480=>x"00015",
481=>x"00015",
482=>x"00014",
483=>x"00014",
484=>x"00014",
485=>x"00014",
486=>x"00014",
487=>x"00014",
488=>x"00014",
489=>x"00014",
490=>x"00014",
491=>x"00014",
492=>x"00014",
493=>x"00014",
494=>x"00014",
495=>x"00014",
496=>x"00014",
497=>x"00014",
498=>x"00014",
499=>x"00014",
500=>x"00014",
501=>x"00014",
502=>x"00014",
503=>x"00014",
504=>x"00014",
505=>x"00014",
506=>x"00014",
507=>x"00014",
508=>x"00014",
509=>x"00014",
510=>x"00014",
511=>x"00014",
512=>x"00014",
513=>x"00013",
514=>x"00013",
515=>x"00013",
516=>x"00013",
517=>x"00013",
518=>x"00013",
519=>x"00013",
520=>x"00013",
521=>x"00013",
522=>x"00013",
523=>x"00013",
524=>x"00013",
525=>x"00013",
526=>x"00013",
527=>x"00013",
528=>x"00013",
529=>x"00013",
530=>x"00013",
531=>x"00013",
532=>x"00013",
533=>x"00013",
534=>x"00013",
535=>x"00013",
536=>x"00013",
537=>x"00013",
538=>x"00013",
539=>x"00013",
540=>x"00013",
541=>x"00013",
542=>x"00013",
543=>x"00013",
544=>x"00013",
545=>x"00013",
546=>x"00012",
547=>x"00012",
548=>x"00012",
549=>x"00012",
550=>x"00012",
551=>x"00012",
552=>x"00012",
553=>x"00012",
554=>x"00012",
555=>x"00012",
556=>x"00012",
557=>x"00012",
558=>x"00012",
559=>x"00012",
560=>x"00012",
561=>x"00012",
562=>x"00012",
563=>x"00012",
564=>x"00012",
565=>x"00012",
566=>x"00012",
567=>x"00012",
568=>x"00012",
569=>x"00012",
570=>x"00012",
571=>x"00012",
572=>x"00012",
573=>x"00012",
574=>x"00012",
575=>x"00012",
576=>x"00012",
577=>x"00012",
578=>x"00012",
579=>x"00012",
580=>x"00012",
581=>x"00012",
582=>x"00012",
583=>x"00012",
584=>x"00011",
585=>x"00011",
586=>x"00011",
587=>x"00011",
588=>x"00011",
589=>x"00011",
590=>x"00011",
591=>x"00011",
592=>x"00011",
593=>x"00011",
594=>x"00011",
595=>x"00011",
596=>x"00011",
597=>x"00011",
598=>x"00011",
599=>x"00011",
600=>x"00011",
601=>x"00011",
602=>x"00011",
603=>x"00011",
604=>x"00011",
605=>x"00011",
606=>x"00011",
607=>x"00011",
608=>x"00011",
609=>x"00011",
610=>x"00011",
611=>x"00011",
612=>x"00011",
613=>x"00011",
614=>x"00011",
615=>x"00011",
616=>x"00011",
617=>x"00011",
618=>x"00011",
619=>x"00011",
620=>x"00011",
621=>x"00011",
622=>x"00011",
623=>x"00011",
624=>x"00011",
625=>x"00010",
626=>x"00010",
627=>x"00010",
628=>x"00010",
629=>x"00010",
630=>x"00010",
631=>x"00010",
632=>x"00010",
633=>x"00010",
634=>x"00010",
635=>x"00010",
636=>x"00010",
637=>x"00010",
638=>x"00010",
639=>x"00010",
640=>x"00010",
641=>x"00010",
642=>x"00010",
643=>x"00010",
644=>x"00010",
645=>x"00010",
646=>x"00010",
647=>x"00010",
648=>x"00010",
649=>x"00010",
650=>x"00010",
651=>x"00010",
652=>x"00010",
653=>x"00010",
654=>x"00010",
655=>x"00010",
656=>x"00010",
657=>x"00010",
658=>x"00010",
659=>x"00010",
660=>x"00010",
661=>x"00010",
662=>x"00010",
663=>x"00010",
664=>x"00010",
665=>x"00010",
666=>x"00010",
667=>x"00010",
668=>x"00010",
669=>x"00010",
670=>x"00010",
671=>x"00010",
672=>x"00010",
673=>x"0000f",
674=>x"0000f",
675=>x"0000f",
676=>x"0000f",
677=>x"0000f",
678=>x"0000f",
679=>x"0000f",
680=>x"0000f",
681=>x"0000f",
682=>x"0000f",
683=>x"0000f",
684=>x"0000f",
685=>x"0000f",
686=>x"0000f",
687=>x"0000f",
688=>x"0000f",
689=>x"0000f",
690=>x"0000f",
691=>x"0000f",
692=>x"0000f",
693=>x"0000f",
694=>x"0000f",
695=>x"0000f",
696=>x"0000f",
697=>x"0000f",
698=>x"0000f",
699=>x"0000f",
700=>x"0000f",
701=>x"0000f",
702=>x"0000f",
703=>x"0000f",
704=>x"0000f",
705=>x"0000f",
706=>x"0000f",
707=>x"0000f",
708=>x"0000f",
709=>x"0000f",
710=>x"0000f",
711=>x"0000f",
712=>x"0000f",
713=>x"0000f",
714=>x"0000f",
715=>x"0000f",
716=>x"0000f",
717=>x"0000f",
718=>x"0000f",
719=>x"0000f",
720=>x"0000f",
721=>x"0000f",
722=>x"0000f",
723=>x"0000f",
724=>x"0000f",
725=>x"0000f",
726=>x"0000e",
727=>x"0000e",
728=>x"0000e",
729=>x"0000e",
730=>x"0000e",
731=>x"0000e",
732=>x"0000e",
733=>x"0000e",
734=>x"0000e",
735=>x"0000e",
736=>x"0000e",
737=>x"0000e",
738=>x"0000e",
739=>x"0000e",
740=>x"0000e",
741=>x"0000e",
742=>x"0000e",
743=>x"0000e",
744=>x"0000e",
745=>x"0000e",
746=>x"0000e",
747=>x"0000e",
748=>x"0000e",
749=>x"0000e",
750=>x"0000e",
751=>x"0000e",
752=>x"0000e",
753=>x"0000e",
754=>x"0000e",
755=>x"0000e",
756=>x"0000e",
757=>x"0000e",
758=>x"0000e",
759=>x"0000e",
760=>x"0000e",
761=>x"0000e",
762=>x"0000e",
763=>x"0000e",
764=>x"0000e",
765=>x"0000e",
766=>x"0000e",
767=>x"0000e",
768=>x"0000e",
769=>x"0000e",
770=>x"0000e",
771=>x"0000e",
772=>x"0000e",
773=>x"0000e",
774=>x"0000e",
775=>x"0000e",
776=>x"0000e",
777=>x"0000e",
778=>x"0000e",
779=>x"0000e",
780=>x"0000e",
781=>x"0000e",
782=>x"0000e",
783=>x"0000e",
784=>x"0000e",
785=>x"0000e",
786=>x"0000e",
787=>x"0000d",
788=>x"0000d",
789=>x"0000d",
790=>x"0000d",
791=>x"0000d",
792=>x"0000d",
793=>x"0000d",
794=>x"0000d",
795=>x"0000d",
796=>x"0000d",
797=>x"0000d",
798=>x"0000d",
799=>x"0000d",
800=>x"0000d",
801=>x"0000d",
802=>x"0000d",
803=>x"0000d",
804=>x"0000d",
805=>x"0000d",
806=>x"0000d",
807=>x"0000d",
808=>x"0000d",
809=>x"0000d",
810=>x"0000d",
811=>x"0000d",
812=>x"0000d",
813=>x"0000d",
814=>x"0000d",
815=>x"0000d",
816=>x"0000d",
817=>x"0000d",
818=>x"0000d",
819=>x"0000d",
820=>x"0000d",
821=>x"0000d",
822=>x"0000d",
823=>x"0000d",
824=>x"0000d",
825=>x"0000d",
826=>x"0000d",
827=>x"0000d",
828=>x"0000d",
829=>x"0000d",
830=>x"0000d",
831=>x"0000d",
832=>x"0000d",
833=>x"0000d",
834=>x"0000d",
835=>x"0000d",
836=>x"0000d",
837=>x"0000d",
838=>x"0000d",
839=>x"0000d",
840=>x"0000d",
841=>x"0000d",
842=>x"0000d",
843=>x"0000d",
844=>x"0000d",
845=>x"0000d",
846=>x"0000d",
847=>x"0000d",
848=>x"0000d",
849=>x"0000d",
850=>x"0000d",
851=>x"0000d",
852=>x"0000d",
853=>x"0000d",
854=>x"0000d",
855=>x"0000d",
856=>x"0000d",
857=>x"0000c",
858=>x"0000c",
859=>x"0000c",
860=>x"0000c",
861=>x"0000c",
862=>x"0000c",
863=>x"0000c",
864=>x"0000c",
865=>x"0000c",
866=>x"0000c",
867=>x"0000c",
868=>x"0000c",
869=>x"0000c",
870=>x"0000c",
871=>x"0000c",
872=>x"0000c",
873=>x"0000c",
874=>x"0000c",
875=>x"0000c",
876=>x"0000c",
877=>x"0000c",
878=>x"0000c",
879=>x"0000c",
880=>x"0000c",
881=>x"0000c",
882=>x"0000c",
883=>x"0000c",
884=>x"0000c",
885=>x"0000c",
886=>x"0000c",
887=>x"0000c",
888=>x"0000c",
889=>x"0000c",
890=>x"0000c",
891=>x"0000c",
892=>x"0000c",
893=>x"0000c",
894=>x"0000c",
895=>x"0000c",
896=>x"0000c",
897=>x"0000c",
898=>x"0000c",
899=>x"0000c",
900=>x"0000c",
901=>x"0000c",
902=>x"0000c",
903=>x"0000c",
904=>x"0000c",
905=>x"0000c",
906=>x"0000c",
907=>x"0000c",
908=>x"0000c",
909=>x"0000c",
910=>x"0000c",
911=>x"0000c",
912=>x"0000c",
913=>x"0000c",
914=>x"0000c",
915=>x"0000c",
916=>x"0000c",
917=>x"0000c",
918=>x"0000c",
919=>x"0000c",
920=>x"0000c",
921=>x"0000c",
922=>x"0000c",
923=>x"0000c",
924=>x"0000c",
925=>x"0000c",
926=>x"0000c",
927=>x"0000c",
928=>x"0000c",
929=>x"0000c",
930=>x"0000c",
931=>x"0000c",
932=>x"0000c",
933=>x"0000c",
934=>x"0000c",
935=>x"0000c",
936=>x"0000c",
937=>x"0000c",
938=>x"0000c",
939=>x"0000b",
940=>x"0000b",
941=>x"0000b",
942=>x"0000b",
943=>x"0000b",
944=>x"0000b",
945=>x"0000b",
946=>x"0000b",
947=>x"0000b",
948=>x"0000b",
949=>x"0000b",
950=>x"0000b",
951=>x"0000b",
952=>x"0000b",
953=>x"0000b",
954=>x"0000b",
955=>x"0000b",
956=>x"0000b",
957=>x"0000b",
958=>x"0000b",
959=>x"0000b",
960=>x"0000b",
961=>x"0000b",
962=>x"0000b",
963=>x"0000b",
964=>x"0000b",
965=>x"0000b",
966=>x"0000b",
967=>x"0000b",
968=>x"0000b",
969=>x"0000b",
970=>x"0000b",
971=>x"0000b",
972=>x"0000b",
973=>x"0000b",
974=>x"0000b",
975=>x"0000b",
976=>x"0000b",
977=>x"0000b",
978=>x"0000b",
979=>x"0000b",
980=>x"0000b",
981=>x"0000b",
982=>x"0000b",
983=>x"0000b",
984=>x"0000b",
985=>x"0000b",
986=>x"0000b",
987=>x"0000b",
988=>x"0000b",
989=>x"0000b",
990=>x"0000b",
991=>x"0000b",
992=>x"0000b",
993=>x"0000b",
994=>x"0000b",
995=>x"0000b",
996=>x"0000b",
997=>x"0000b",
998=>x"0000b",
999=>x"0000b",
1000=>x"0000b",
1001=>x"0000b",
1002=>x"0000b",
1003=>x"0000b",
1004=>x"0000b",
1005=>x"0000b",
1006=>x"0000b",
1007=>x"0000b",
1008=>x"0000b",
1009=>x"0000b",
1010=>x"0000b",
1011=>x"0000b",
1012=>x"0000b",
1013=>x"0000b",
1014=>x"0000b",
1015=>x"0000b",
1016=>x"0000b",
1017=>x"0000b",
1018=>x"0000b",
1019=>x"0000b",
1020=>x"0000b",
1021=>x"0000b",
1022=>x"0000b",
1023=>x"0000b",
1024=>x"0000b",
1025=>x"0000b",
1026=>x"0000b",
1027=>x"0000b",
1028=>x"0000b",
1029=>x"0000b",
1030=>x"0000b",
1031=>x"0000b",
1032=>x"0000b",
1033=>x"0000b",
1034=>x"0000b",
1035=>x"0000b",
1036=>x"0000a",
1037=>x"0000a",
1038=>x"0000a",
1039=>x"0000a",
1040=>x"0000a",
1041=>x"0000a",
1042=>x"0000a",
1043=>x"0000a",
1044=>x"0000a",
1045=>x"0000a",
1046=>x"0000a",
1047=>x"0000a",
1048=>x"0000a",
1049=>x"0000a",
1050=>x"0000a",
1051=>x"0000a",
1052=>x"0000a",
1053=>x"0000a",
1054=>x"0000a",
1055=>x"0000a",
1056=>x"0000a",
1057=>x"0000a",
1058=>x"0000a",
1059=>x"0000a",
1060=>x"0000a",
1061=>x"0000a",
1062=>x"0000a",
1063=>x"0000a",
1064=>x"0000a",
1065=>x"0000a",
1066=>x"0000a",
1067=>x"0000a",
1068=>x"0000a",
1069=>x"0000a",
1070=>x"0000a",
1071=>x"0000a",
1072=>x"0000a",
1073=>x"0000a",
1074=>x"0000a",
1075=>x"0000a",
1076=>x"0000a",
1077=>x"0000a",
1078=>x"0000a",
1079=>x"0000a",
1080=>x"0000a",
1081=>x"0000a",
1082=>x"0000a",
1083=>x"0000a",
1084=>x"0000a",
1085=>x"0000a",
1086=>x"0000a",
1087=>x"0000a",
1088=>x"0000a",
1089=>x"0000a",
1090=>x"0000a",
1091=>x"0000a",
1092=>x"0000a",
1093=>x"0000a",
1094=>x"0000a",
1095=>x"0000a",
1096=>x"0000a",
1097=>x"0000a",
1098=>x"0000a",
1099=>x"0000a",
1100=>x"0000a",
1101=>x"0000a",
1102=>x"0000a",
1103=>x"0000a",
1104=>x"0000a",
1105=>x"0000a",
1106=>x"0000a",
1107=>x"0000a",
1108=>x"0000a",
1109=>x"0000a",
1110=>x"0000a",
1111=>x"0000a",
1112=>x"0000a",
1113=>x"0000a",
1114=>x"0000a",
1115=>x"0000a",
1116=>x"0000a",
1117=>x"0000a",
1118=>x"0000a",
1119=>x"0000a",
1120=>x"0000a",
1121=>x"0000a",
1122=>x"0000a",
1123=>x"0000a",
1124=>x"0000a",
1125=>x"0000a",
1126=>x"0000a",
1127=>x"0000a",
1128=>x"0000a",
1129=>x"0000a",
1130=>x"0000a",
1131=>x"0000a",
1132=>x"0000a",
1133=>x"0000a",
1134=>x"0000a",
1135=>x"0000a",
1136=>x"0000a",
1137=>x"0000a",
1138=>x"0000a",
1139=>x"0000a",
1140=>x"0000a",
1141=>x"0000a",
1142=>x"0000a",
1143=>x"0000a",
1144=>x"0000a",
1145=>x"0000a",
1146=>x"0000a",
1147=>x"0000a",
1148=>x"0000a",
1149=>x"0000a",
1150=>x"0000a",
1151=>x"0000a",
1152=>x"0000a",
1153=>x"00009",
1154=>x"00009",
1155=>x"00009",
1156=>x"00009",
1157=>x"00009",
1158=>x"00009",
1159=>x"00009",
1160=>x"00009",
1161=>x"00009",
1162=>x"00009",
1163=>x"00009",
1164=>x"00009",
1165=>x"00009",
1166=>x"00009",
1167=>x"00009",
1168=>x"00009",
1169=>x"00009",
1170=>x"00009",
1171=>x"00009",
1172=>x"00009",
1173=>x"00009",
1174=>x"00009",
1175=>x"00009",
1176=>x"00009",
1177=>x"00009",
1178=>x"00009",
1179=>x"00009",
1180=>x"00009",
1181=>x"00009",
1182=>x"00009",
1183=>x"00009",
1184=>x"00009",
1185=>x"00009",
1186=>x"00009",
1187=>x"00009",
1188=>x"00009",
1189=>x"00009",
1190=>x"00009",
1191=>x"00009",
1192=>x"00009",
1193=>x"00009",
1194=>x"00009",
1195=>x"00009",
1196=>x"00009",
1197=>x"00009",
1198=>x"00009",
1199=>x"00009",
1200=>x"00009",
1201=>x"00009",
1202=>x"00009",
1203=>x"00009",
1204=>x"00009",
1205=>x"00009",
1206=>x"00009",
1207=>x"00009",
1208=>x"00009",
1209=>x"00009",
1210=>x"00009",
1211=>x"00009",
1212=>x"00009",
1213=>x"00009",
1214=>x"00009",
1215=>x"00009",
1216=>x"00009",
1217=>x"00009",
1218=>x"00009",
1219=>x"00009",
1220=>x"00009",
1221=>x"00009",
1222=>x"00009",
1223=>x"00009",
1224=>x"00009",
1225=>x"00009",
1226=>x"00009",
1227=>x"00009",
1228=>x"00009",
1229=>x"00009",
1230=>x"00009",
1231=>x"00009",
1232=>x"00009",
1233=>x"00009",
1234=>x"00009",
1235=>x"00009",
1236=>x"00009",
1237=>x"00009",
1238=>x"00009",
1239=>x"00009",
1240=>x"00009",
1241=>x"00009",
1242=>x"00009",
1243=>x"00009",
1244=>x"00009",
1245=>x"00009",
1246=>x"00009",
1247=>x"00009",
1248=>x"00009",
1249=>x"00009",
1250=>x"00009",
1251=>x"00009",
1252=>x"00009",
1253=>x"00009",
1254=>x"00009",
1255=>x"00009",
1256=>x"00009",
1257=>x"00009",
1258=>x"00009",
1259=>x"00009",
1260=>x"00009",
1261=>x"00009",
1262=>x"00009",
1263=>x"00009",
1264=>x"00009",
1265=>x"00009",
1266=>x"00009",
1267=>x"00009",
1268=>x"00009",
1269=>x"00009",
1270=>x"00009",
1271=>x"00009",
1272=>x"00009",
1273=>x"00009",
1274=>x"00009",
1275=>x"00009",
1276=>x"00009",
1277=>x"00009",
1278=>x"00009",
1279=>x"00009",
1280=>x"00009",
1281=>x"00009",
1282=>x"00009",
1283=>x"00009",
1284=>x"00009",
1285=>x"00009",
1286=>x"00009",
1287=>x"00009",
1288=>x"00009",
1289=>x"00009",
1290=>x"00009",
1291=>x"00009",
1292=>x"00009",
1293=>x"00009",
1294=>x"00009",
1295=>x"00008",
1296=>x"00008",
1297=>x"00008",
1298=>x"00008",
1299=>x"00008",
1300=>x"00008",
1301=>x"00008",
1302=>x"00008",
1303=>x"00008",
1304=>x"00008",
1305=>x"00008",
1306=>x"00008",
1307=>x"00008",
1308=>x"00008",
1309=>x"00008",
1310=>x"00008",
1311=>x"00008",
1312=>x"00008",
1313=>x"00008",
1314=>x"00008",
1315=>x"00008",
1316=>x"00008",
1317=>x"00008",
1318=>x"00008",
1319=>x"00008",
1320=>x"00008",
1321=>x"00008",
1322=>x"00008",
1323=>x"00008",
1324=>x"00008",
1325=>x"00008",
1326=>x"00008",
1327=>x"00008",
1328=>x"00008",
1329=>x"00008",
1330=>x"00008",
1331=>x"00008",
1332=>x"00008",
1333=>x"00008",
1334=>x"00008",
1335=>x"00008",
1336=>x"00008",
1337=>x"00008",
1338=>x"00008",
1339=>x"00008",
1340=>x"00008",
1341=>x"00008",
1342=>x"00008",
1343=>x"00008",
1344=>x"00008",
1345=>x"00008",
1346=>x"00008",
1347=>x"00008",
1348=>x"00008",
1349=>x"00008",
1350=>x"00008",
1351=>x"00008",
1352=>x"00008",
1353=>x"00008",
1354=>x"00008",
1355=>x"00008",
1356=>x"00008",
1357=>x"00008",
1358=>x"00008",
1359=>x"00008",
1360=>x"00008",
1361=>x"00008",
1362=>x"00008",
1363=>x"00008",
1364=>x"00008",
1365=>x"00008",
1366=>x"00008",
1367=>x"00008",
1368=>x"00008",
1369=>x"00008",
1370=>x"00008",
1371=>x"00008",
1372=>x"00008",
1373=>x"00008",
1374=>x"00008",
1375=>x"00008",
1376=>x"00008",
1377=>x"00008",
1378=>x"00008",
1379=>x"00008",
1380=>x"00008",
1381=>x"00008",
1382=>x"00008",
1383=>x"00008",
1384=>x"00008",
1385=>x"00008",
1386=>x"00008",
1387=>x"00008",
1388=>x"00008",
1389=>x"00008",
1390=>x"00008",
1391=>x"00008",
1392=>x"00008",
1393=>x"00008",
1394=>x"00008",
1395=>x"00008",
1396=>x"00008",
1397=>x"00008",
1398=>x"00008",
1399=>x"00008",
1400=>x"00008",
1401=>x"00008",
1402=>x"00008",
1403=>x"00008",
1404=>x"00008",
1405=>x"00008",
1406=>x"00008",
1407=>x"00008",
1408=>x"00008",
1409=>x"00008",
1410=>x"00008",
1411=>x"00008",
1412=>x"00008",
1413=>x"00008",
1414=>x"00008",
1415=>x"00008",
1416=>x"00008",
1417=>x"00008",
1418=>x"00008",
1419=>x"00008",
1420=>x"00008",
1421=>x"00008",
1422=>x"00008",
1423=>x"00008",
1424=>x"00008",
1425=>x"00008",
1426=>x"00008",
1427=>x"00008",
1428=>x"00008",
1429=>x"00008",
1430=>x"00008",
1431=>x"00008",
1432=>x"00008",
1433=>x"00008",
1434=>x"00008",
1435=>x"00008",
1436=>x"00008",
1437=>x"00008",
1438=>x"00008",
1439=>x"00008",
1440=>x"00008",
1441=>x"00008",
1442=>x"00008",
1443=>x"00008",
1444=>x"00008",
1445=>x"00008",
1446=>x"00008",
1447=>x"00008",
1448=>x"00008",
1449=>x"00008",
1450=>x"00008",
1451=>x"00008",
1452=>x"00008",
1453=>x"00008",
1454=>x"00008",
1455=>x"00008",
1456=>x"00008",
1457=>x"00008",
1458=>x"00008",
1459=>x"00008",
1460=>x"00008",
1461=>x"00008",
1462=>x"00008",
1463=>x"00008",
1464=>x"00008",
1465=>x"00008",
1466=>x"00008",
1467=>x"00008",
1468=>x"00008",
1469=>x"00008",
1470=>x"00008",
1471=>x"00008",
1472=>x"00008",
1473=>x"00007",
1474=>x"00007",
1475=>x"00007",
1476=>x"00007",
1477=>x"00007",
1478=>x"00007",
1479=>x"00007",
1480=>x"00007",
1481=>x"00007",
1482=>x"00007",
1483=>x"00007",
1484=>x"00007",
1485=>x"00007",
1486=>x"00007",
1487=>x"00007",
1488=>x"00007",
1489=>x"00007",
1490=>x"00007",
1491=>x"00007",
1492=>x"00007",
1493=>x"00007",
1494=>x"00007",
1495=>x"00007",
1496=>x"00007",
1497=>x"00007",
1498=>x"00007",
1499=>x"00007",
1500=>x"00007",
1501=>x"00007",
1502=>x"00007",
1503=>x"00007",
1504=>x"00007",
1505=>x"00007",
1506=>x"00007",
1507=>x"00007",
1508=>x"00007",
1509=>x"00007",
1510=>x"00007",
1511=>x"00007",
1512=>x"00007",
1513=>x"00007",
1514=>x"00007",
1515=>x"00007",
1516=>x"00007",
1517=>x"00007",
1518=>x"00007",
1519=>x"00007",
1520=>x"00007",
1521=>x"00007",
1522=>x"00007",
1523=>x"00007",
1524=>x"00007",
1525=>x"00007",
1526=>x"00007",
1527=>x"00007",
1528=>x"00007",
1529=>x"00007",
1530=>x"00007",
1531=>x"00007",
1532=>x"00007",
1533=>x"00007",
1534=>x"00007",
1535=>x"00007",
1536=>x"00007",
1537=>x"00007",
1538=>x"00007",
1539=>x"00007",
1540=>x"00007",
1541=>x"00007",
1542=>x"00007",
1543=>x"00007",
1544=>x"00007",
1545=>x"00007",
1546=>x"00007",
1547=>x"00007",
1548=>x"00007",
1549=>x"00007",
1550=>x"00007",
1551=>x"00007",
1552=>x"00007",
1553=>x"00007",
1554=>x"00007",
1555=>x"00007",
1556=>x"00007",
1557=>x"00007",
1558=>x"00007",
1559=>x"00007",
1560=>x"00007",
1561=>x"00007",
1562=>x"00007",
1563=>x"00007",
1564=>x"00007",
1565=>x"00007",
1566=>x"00007",
1567=>x"00007",
1568=>x"00007",
1569=>x"00007",
1570=>x"00007",
1571=>x"00007",
1572=>x"00007",
1573=>x"00007",
1574=>x"00007",
1575=>x"00007",
1576=>x"00007",
1577=>x"00007",
1578=>x"00007",
1579=>x"00007",
1580=>x"00007",
1581=>x"00007",
1582=>x"00007",
1583=>x"00007",
1584=>x"00007",
1585=>x"00007",
1586=>x"00007",
1587=>x"00007",
1588=>x"00007",
1589=>x"00007",
1590=>x"00007",
1591=>x"00007",
1592=>x"00007",
1593=>x"00007",
1594=>x"00007",
1595=>x"00007",
1596=>x"00007",
1597=>x"00007",
1598=>x"00007",
1599=>x"00007",
1600=>x"00007",
1601=>x"00007",
1602=>x"00007",
1603=>x"00007",
1604=>x"00007",
1605=>x"00007",
1606=>x"00007",
1607=>x"00007",
1608=>x"00007",
1609=>x"00007",
1610=>x"00007",
1611=>x"00007",
1612=>x"00007",
1613=>x"00007",
1614=>x"00007",
1615=>x"00007",
1616=>x"00007",
1617=>x"00007",
1618=>x"00007",
1619=>x"00007",
1620=>x"00007",
1621=>x"00007",
1622=>x"00007",
1623=>x"00007",
1624=>x"00007",
1625=>x"00007",
1626=>x"00007",
1627=>x"00007",
1628=>x"00007",
1629=>x"00007",
1630=>x"00007",
1631=>x"00007",
1632=>x"00007",
1633=>x"00007",
1634=>x"00007",
1635=>x"00007",
1636=>x"00007",
1637=>x"00007",
1638=>x"00007",
1639=>x"00007",
1640=>x"00007",
1641=>x"00007",
1642=>x"00007",
1643=>x"00007",
1644=>x"00007",
1645=>x"00007",
1646=>x"00007",
1647=>x"00007",
1648=>x"00007",
1649=>x"00007",
1650=>x"00007",
1651=>x"00007",
1652=>x"00007",
1653=>x"00007",
1654=>x"00007",
1655=>x"00007",
1656=>x"00007",
1657=>x"00007",
1658=>x"00007",
1659=>x"00007",
1660=>x"00007",
1661=>x"00007",
1662=>x"00007",
1663=>x"00007",
1664=>x"00007",
1665=>x"00007",
1666=>x"00007",
1667=>x"00007",
1668=>x"00007",
1669=>x"00007",
1670=>x"00007",
1671=>x"00007",
1672=>x"00007",
1673=>x"00007",
1674=>x"00007",
1675=>x"00007",
1676=>x"00007",
1677=>x"00007",
1678=>x"00007",
1679=>x"00007",
1680=>x"00007",
1681=>x"00007",
1682=>x"00007",
1683=>x"00007",
1684=>x"00007",
1685=>x"00007",
1686=>x"00007",
1687=>x"00007",
1688=>x"00007",
1689=>x"00007",
1690=>x"00007",
1691=>x"00007",
1692=>x"00007",
1693=>x"00007",
1694=>x"00007",
1695=>x"00007",
1696=>x"00007",
1697=>x"00007",
1698=>x"00007",
1699=>x"00007",
1700=>x"00007",
1701=>x"00006",
1702=>x"00006",
1703=>x"00006",
1704=>x"00006",
1705=>x"00006",
1706=>x"00006",
1707=>x"00006",
1708=>x"00006",
1709=>x"00006",
1710=>x"00006",
1711=>x"00006",
1712=>x"00006",
1713=>x"00006",
1714=>x"00006",
1715=>x"00006",
1716=>x"00006",
1717=>x"00006",
1718=>x"00006",
1719=>x"00006",
1720=>x"00006",
1721=>x"00006",
1722=>x"00006",
1723=>x"00006",
1724=>x"00006",
1725=>x"00006",
1726=>x"00006",
1727=>x"00006",
1728=>x"00006",
1729=>x"00006",
1730=>x"00006",
1731=>x"00006",
1732=>x"00006",
1733=>x"00006",
1734=>x"00006",
1735=>x"00006",
1736=>x"00006",
1737=>x"00006",
1738=>x"00006",
1739=>x"00006",
1740=>x"00006",
1741=>x"00006",
1742=>x"00006",
1743=>x"00006",
1744=>x"00006",
1745=>x"00006",
1746=>x"00006",
1747=>x"00006",
1748=>x"00006",
1749=>x"00006",
1750=>x"00006",
1751=>x"00006",
1752=>x"00006",
1753=>x"00006",
1754=>x"00006",
1755=>x"00006",
1756=>x"00006",
1757=>x"00006",
1758=>x"00006",
1759=>x"00006",
1760=>x"00006",
1761=>x"00006",
1762=>x"00006",
1763=>x"00006",
1764=>x"00006",
1765=>x"00006",
1766=>x"00006",
1767=>x"00006",
1768=>x"00006",
1769=>x"00006",
1770=>x"00006",
1771=>x"00006",
1772=>x"00006",
1773=>x"00006",
1774=>x"00006",
1775=>x"00006",
1776=>x"00006",
1777=>x"00006",
1778=>x"00006",
1779=>x"00006",
1780=>x"00006",
1781=>x"00006",
1782=>x"00006",
1783=>x"00006",
1784=>x"00006",
1785=>x"00006",
1786=>x"00006",
1787=>x"00006",
1788=>x"00006",
1789=>x"00006",
1790=>x"00006",
1791=>x"00006",
1792=>x"00006",
1793=>x"00006",
1794=>x"00006",
1795=>x"00006",
1796=>x"00006",
1797=>x"00006",
1798=>x"00006",
1799=>x"00006",
1800=>x"00006",
1801=>x"00006",
1802=>x"00006",
1803=>x"00006",
1804=>x"00006",
1805=>x"00006",
1806=>x"00006",
1807=>x"00006",
1808=>x"00006",
1809=>x"00006",
1810=>x"00006",
1811=>x"00006",
1812=>x"00006",
1813=>x"00006",
1814=>x"00006",
1815=>x"00006",
1816=>x"00006",
1817=>x"00006",
1818=>x"00006",
1819=>x"00006",
1820=>x"00006",
1821=>x"00006",
1822=>x"00006",
1823=>x"00006",
1824=>x"00006",
1825=>x"00006",
1826=>x"00006",
1827=>x"00006",
1828=>x"00006",
1829=>x"00006",
1830=>x"00006",
1831=>x"00006",
1832=>x"00006",
1833=>x"00006",
1834=>x"00006",
1835=>x"00006",
1836=>x"00006",
1837=>x"00006",
1838=>x"00006",
1839=>x"00006",
1840=>x"00006",
1841=>x"00006",
1842=>x"00006",
1843=>x"00006",
1844=>x"00006",
1845=>x"00006",
1846=>x"00006",
1847=>x"00006",
1848=>x"00006",
1849=>x"00006",
1850=>x"00006",
1851=>x"00006",
1852=>x"00006",
1853=>x"00006",
1854=>x"00006",
1855=>x"00006",
1856=>x"00006",
1857=>x"00006",
1858=>x"00006",
1859=>x"00006",
1860=>x"00006",
1861=>x"00006",
1862=>x"00006",
1863=>x"00006",
1864=>x"00006",
1865=>x"00006",
1866=>x"00006",
1867=>x"00006",
1868=>x"00006",
1869=>x"00006",
1870=>x"00006",
1871=>x"00006",
1872=>x"00006",
1873=>x"00006",
1874=>x"00006",
1875=>x"00006",
1876=>x"00006",
1877=>x"00006",
1878=>x"00006",
1879=>x"00006",
1880=>x"00006",
1881=>x"00006",
1882=>x"00006",
1883=>x"00006",
1884=>x"00006",
1885=>x"00006",
1886=>x"00006",
1887=>x"00006",
1888=>x"00006",
1889=>x"00006",
1890=>x"00006",
1891=>x"00006",
1892=>x"00006",
1893=>x"00006",
1894=>x"00006",
1895=>x"00006",
1896=>x"00006",
1897=>x"00006",
1898=>x"00006",
1899=>x"00006",
1900=>x"00006",
1901=>x"00006",
1902=>x"00006",
1903=>x"00006",
1904=>x"00006",
1905=>x"00006",
1906=>x"00006",
1907=>x"00006",
1908=>x"00006",
1909=>x"00006",
1910=>x"00006",
1911=>x"00006",
1912=>x"00006",
1913=>x"00006",
1914=>x"00006",
1915=>x"00006",
1916=>x"00006",
1917=>x"00006",
1918=>x"00006",
1919=>x"00006",
1920=>x"00006",
1921=>x"00006",
1922=>x"00006",
1923=>x"00006",
1924=>x"00006",
1925=>x"00006",
1926=>x"00006",
1927=>x"00006",
1928=>x"00006",
1929=>x"00006",
1930=>x"00006",
1931=>x"00006",
1932=>x"00006",
1933=>x"00006",
1934=>x"00006",
1935=>x"00006",
1936=>x"00006",
1937=>x"00006",
1938=>x"00006",
1939=>x"00006",
1940=>x"00006",
1941=>x"00006",
1942=>x"00006",
1943=>x"00006",
1944=>x"00006",
1945=>x"00006",
1946=>x"00006",
1947=>x"00006",
1948=>x"00006",
1949=>x"00006",
1950=>x"00006",
1951=>x"00006",
1952=>x"00006",
1953=>x"00006",
1954=>x"00006",
1955=>x"00006",
1956=>x"00006",
1957=>x"00006",
1958=>x"00006",
1959=>x"00006",
1960=>x"00006",
1961=>x"00006",
1962=>x"00006",
1963=>x"00006",
1964=>x"00006",
1965=>x"00006",
1966=>x"00006",
1967=>x"00006",
1968=>x"00006",
1969=>x"00006",
1970=>x"00006",
1971=>x"00006",
1972=>x"00006",
1973=>x"00006",
1974=>x"00006",
1975=>x"00006",
1976=>x"00006",
1977=>x"00006",
1978=>x"00006",
1979=>x"00006",
1980=>x"00006",
1981=>x"00006",
1982=>x"00006",
1983=>x"00006",
1984=>x"00006",
1985=>x"00006",
1986=>x"00006",
1987=>x"00006",
1988=>x"00006",
1989=>x"00006",
1990=>x"00006",
1991=>x"00006",
1992=>x"00006",
1993=>x"00006",
1994=>x"00006",
1995=>x"00006",
1996=>x"00006",
1997=>x"00006",
1998=>x"00006",
1999=>x"00006",
2000=>x"00006",
2001=>x"00006",
2002=>x"00006",
2003=>x"00006",
2004=>x"00006",
2005=>x"00006",
2006=>x"00005",
2007=>x"00005",
2008=>x"00005",
2009=>x"00005",
2010=>x"00005",
2011=>x"00005",
2012=>x"00005",
2013=>x"00005",
2014=>x"00005",
2015=>x"00005",
2016=>x"00005",
2017=>x"00005",
2018=>x"00005",
2019=>x"00005",
2020=>x"00005",
2021=>x"00005",
2022=>x"00005",
2023=>x"00005",
2024=>x"00005",
2025=>x"00005",
2026=>x"00005",
2027=>x"00005",
2028=>x"00005",
2029=>x"00005",
2030=>x"00005",
2031=>x"00005",
2032=>x"00005",
2033=>x"00005",
2034=>x"00005",
2035=>x"00005",
2036=>x"00005",
2037=>x"00005",
2038=>x"00005",
2039=>x"00005",
2040=>x"00005",
2041=>x"00005",
2042=>x"00005",
2043=>x"00005",
2044=>x"00005",
2045=>x"00005",
2046=>x"00005",
2047=>x"00005",
2048=>x"00005",
2049=>x"00005",
2050=>x"00005",
2051=>x"00005",
2052=>x"00005",
2053=>x"00005",
2054=>x"00005",
2055=>x"00005",
2056=>x"00005",
2057=>x"00005",
2058=>x"00005",
2059=>x"00005",
2060=>x"00005",
2061=>x"00005",
2062=>x"00005",
2063=>x"00005",
2064=>x"00005",
2065=>x"00005",
2066=>x"00005",
2067=>x"00005",
2068=>x"00005",
2069=>x"00005",
2070=>x"00005",
2071=>x"00005",
2072=>x"00005",
2073=>x"00005",
2074=>x"00005",
2075=>x"00005",
2076=>x"00005",
2077=>x"00005",
2078=>x"00005",
2079=>x"00005",
2080=>x"00005",
2081=>x"00005",
2082=>x"00005",
2083=>x"00005",
2084=>x"00005",
2085=>x"00005",
2086=>x"00005",
2087=>x"00005",
2088=>x"00005",
2089=>x"00005",
2090=>x"00005",
2091=>x"00005",
2092=>x"00005",
2093=>x"00005",
2094=>x"00005",
2095=>x"00005",
2096=>x"00005",
2097=>x"00005",
2098=>x"00005",
2099=>x"00005",
2100=>x"00005",
2101=>x"00005",
2102=>x"00005",
2103=>x"00005",
2104=>x"00005",
2105=>x"00005",
2106=>x"00005",
2107=>x"00005",
2108=>x"00005",
2109=>x"00005",
2110=>x"00005",
2111=>x"00005",
2112=>x"00005",
2113=>x"00005",
2114=>x"00005",
2115=>x"00005",
2116=>x"00005",
2117=>x"00005",
2118=>x"00005",
2119=>x"00005",
2120=>x"00005",
2121=>x"00005",
2122=>x"00005",
2123=>x"00005",
2124=>x"00005",
2125=>x"00005",
2126=>x"00005",
2127=>x"00005",
2128=>x"00005",
2129=>x"00005",
2130=>x"00005",
2131=>x"00005",
2132=>x"00005",
2133=>x"00005",
2134=>x"00005",
2135=>x"00005",
2136=>x"00005",
2137=>x"00005",
2138=>x"00005",
2139=>x"00005",
2140=>x"00005",
2141=>x"00005",
2142=>x"00005",
2143=>x"00005",
2144=>x"00005",
2145=>x"00005",
2146=>x"00005",
2147=>x"00005",
2148=>x"00005",
2149=>x"00005",
2150=>x"00005",
2151=>x"00005",
2152=>x"00005",
2153=>x"00005",
2154=>x"00005",
2155=>x"00005",
2156=>x"00005",
2157=>x"00005",
2158=>x"00005",
2159=>x"00005",
2160=>x"00005",
2161=>x"00005",
2162=>x"00005",
2163=>x"00005",
2164=>x"00005",
2165=>x"00005",
2166=>x"00005",
2167=>x"00005",
2168=>x"00005",
2169=>x"00005",
2170=>x"00005",
2171=>x"00005",
2172=>x"00005",
2173=>x"00005",
2174=>x"00005",
2175=>x"00005",
2176=>x"00005",
2177=>x"00005",
2178=>x"00005",
2179=>x"00005",
2180=>x"00005",
2181=>x"00005",
2182=>x"00005",
2183=>x"00005",
2184=>x"00005",
2185=>x"00005",
2186=>x"00005",
2187=>x"00005",
2188=>x"00005",
2189=>x"00005",
2190=>x"00005",
2191=>x"00005",
2192=>x"00005",
2193=>x"00005",
2194=>x"00005",
2195=>x"00005",
2196=>x"00005",
2197=>x"00005",
2198=>x"00005",
2199=>x"00005",
2200=>x"00005",
2201=>x"00005",
2202=>x"00005",
2203=>x"00005",
2204=>x"00005",
2205=>x"00005",
2206=>x"00005",
2207=>x"00005",
2208=>x"00005",
2209=>x"00005",
2210=>x"00005",
2211=>x"00005",
2212=>x"00005",
2213=>x"00005",
2214=>x"00005",
2215=>x"00005",
2216=>x"00005",
2217=>x"00005",
2218=>x"00005",
2219=>x"00005",
2220=>x"00005",
2221=>x"00005",
2222=>x"00005",
2223=>x"00005",
2224=>x"00005",
2225=>x"00005",
2226=>x"00005",
2227=>x"00005",
2228=>x"00005",
2229=>x"00005",
2230=>x"00005",
2231=>x"00005",
2232=>x"00005",
2233=>x"00005",
2234=>x"00005",
2235=>x"00005",
2236=>x"00005",
2237=>x"00005",
2238=>x"00005",
2239=>x"00005",
2240=>x"00005",
2241=>x"00005",
2242=>x"00005",
2243=>x"00005",
2244=>x"00005",
2245=>x"00005",
2246=>x"00005",
2247=>x"00005",
2248=>x"00005",
2249=>x"00005",
2250=>x"00005",
2251=>x"00005",
2252=>x"00005",
2253=>x"00005",
2254=>x"00005",
2255=>x"00005",
2256=>x"00005",
2257=>x"00005",
2258=>x"00005",
2259=>x"00005",
2260=>x"00005",
2261=>x"00005",
2262=>x"00005",
2263=>x"00005",
2264=>x"00005",
2265=>x"00005",
2266=>x"00005",
2267=>x"00005",
2268=>x"00005",
2269=>x"00005",
2270=>x"00005",
2271=>x"00005",
2272=>x"00005",
2273=>x"00005",
2274=>x"00005",
2275=>x"00005",
2276=>x"00005",
2277=>x"00005",
2278=>x"00005",
2279=>x"00005",
2280=>x"00005",
2281=>x"00005",
2282=>x"00005",
2283=>x"00005",
2284=>x"00005",
2285=>x"00005",
2286=>x"00005",
2287=>x"00005",
2288=>x"00005",
2289=>x"00005",
2290=>x"00005",
2291=>x"00005",
2292=>x"00005",
2293=>x"00005",
2294=>x"00005",
2295=>x"00005",
2296=>x"00005",
2297=>x"00005",
2298=>x"00005",
2299=>x"00005",
2300=>x"00005",
2301=>x"00005",
2302=>x"00005",
2303=>x"00005",
2304=>x"00005",
2305=>x"00005",
2306=>x"00005",
2307=>x"00005",
2308=>x"00005",
2309=>x"00005",
2310=>x"00005",
2311=>x"00005",
2312=>x"00005",
2313=>x"00005",
2314=>x"00005",
2315=>x"00005",
2316=>x"00005",
2317=>x"00005",
2318=>x"00005",
2319=>x"00005",
2320=>x"00005",
2321=>x"00005",
2322=>x"00005",
2323=>x"00005",
2324=>x"00005",
2325=>x"00005",
2326=>x"00005",
2327=>x"00005",
2328=>x"00005",
2329=>x"00005",
2330=>x"00005",
2331=>x"00005",
2332=>x"00005",
2333=>x"00005",
2334=>x"00005",
2335=>x"00005",
2336=>x"00005",
2337=>x"00005",
2338=>x"00005",
2339=>x"00005",
2340=>x"00005",
2341=>x"00005",
2342=>x"00005",
2343=>x"00005",
2344=>x"00005",
2345=>x"00005",
2346=>x"00005",
2347=>x"00005",
2348=>x"00005",
2349=>x"00005",
2350=>x"00005",
2351=>x"00005",
2352=>x"00005",
2353=>x"00005",
2354=>x"00005",
2355=>x"00005",
2356=>x"00005",
2357=>x"00005",
2358=>x"00005",
2359=>x"00005",
2360=>x"00005",
2361=>x"00005",
2362=>x"00005",
2363=>x"00005",
2364=>x"00005",
2365=>x"00005",
2366=>x"00005",
2367=>x"00005",
2368=>x"00005",
2369=>x"00005",
2370=>x"00005",
2371=>x"00005",
2372=>x"00005",
2373=>x"00005",
2374=>x"00005",
2375=>x"00005",
2376=>x"00005",
2377=>x"00005",
2378=>x"00005",
2379=>x"00005",
2380=>x"00005",
2381=>x"00005",
2382=>x"00005",
2383=>x"00005",
2384=>x"00005",
2385=>x"00005",
2386=>x"00005",
2387=>x"00005",
2388=>x"00005",
2389=>x"00005",
2390=>x"00005",
2391=>x"00005",
2392=>x"00005",
2393=>x"00005",
2394=>x"00005",
2395=>x"00005",
2396=>x"00005",
2397=>x"00005",
2398=>x"00005",
2399=>x"00005",
2400=>x"00005",
2401=>x"00005",
2402=>x"00005",
2403=>x"00005",
2404=>x"00005",
2405=>x"00005",
2406=>x"00005",
2407=>x"00005",
2408=>x"00005",
2409=>x"00005",
2410=>x"00005",
2411=>x"00005",
2412=>x"00005",
2413=>x"00005",
2414=>x"00005",
2415=>x"00005",
2416=>x"00005",
2417=>x"00005",
2418=>x"00005",
2419=>x"00005",
2420=>x"00005",
2421=>x"00005",
2422=>x"00005",
2423=>x"00005",
2424=>x"00005",
2425=>x"00005",
2426=>x"00005",
2427=>x"00005",
2428=>x"00005",
2429=>x"00005",
2430=>x"00005",
2431=>x"00005",
2432=>x"00005",
2433=>x"00004",
2434=>x"00004",
2435=>x"00004",
2436=>x"00004",
2437=>x"00004",
2438=>x"00004",
2439=>x"00004",
2440=>x"00004",
2441=>x"00004",
2442=>x"00004",
2443=>x"00004",
2444=>x"00004",
2445=>x"00004",
2446=>x"00004",
2447=>x"00004",
2448=>x"00004",
2449=>x"00004",
2450=>x"00004",
2451=>x"00004",
2452=>x"00004",
2453=>x"00004",
2454=>x"00004",
2455=>x"00004",
2456=>x"00004",
2457=>x"00004",
2458=>x"00004",
2459=>x"00004",
2460=>x"00004",
2461=>x"00004",
2462=>x"00004",
2463=>x"00004",
2464=>x"00004",
2465=>x"00004",
2466=>x"00004",
2467=>x"00004",
2468=>x"00004",
2469=>x"00004",
2470=>x"00004",
2471=>x"00004",
2472=>x"00004",
2473=>x"00004",
2474=>x"00004",
2475=>x"00004",
2476=>x"00004",
2477=>x"00004",
2478=>x"00004",
2479=>x"00004",
2480=>x"00004",
2481=>x"00004",
2482=>x"00004",
2483=>x"00004",
2484=>x"00004",
2485=>x"00004",
2486=>x"00004",
2487=>x"00004",
2488=>x"00004",
2489=>x"00004",
2490=>x"00004",
2491=>x"00004",
2492=>x"00004",
2493=>x"00004",
2494=>x"00004",
2495=>x"00004",
2496=>x"00004",
2497=>x"00004",
2498=>x"00004",
2499=>x"00004",
2500=>x"00004",
2501=>x"00004",
2502=>x"00004",
2503=>x"00004",
2504=>x"00004",
2505=>x"00004",
2506=>x"00004",
2507=>x"00004",
2508=>x"00004",
2509=>x"00004",
2510=>x"00004",
2511=>x"00004",
2512=>x"00004",
2513=>x"00004",
2514=>x"00004",
2515=>x"00004",
2516=>x"00004",
2517=>x"00004",
2518=>x"00004",
2519=>x"00004",
2520=>x"00004",
2521=>x"00004",
2522=>x"00004",
2523=>x"00004",
2524=>x"00004",
2525=>x"00004",
2526=>x"00004",
2527=>x"00004",
2528=>x"00004",
2529=>x"00004",
2530=>x"00004",
2531=>x"00004",
2532=>x"00004",
2533=>x"00004",
2534=>x"00004",
2535=>x"00004",
2536=>x"00004",
2537=>x"00004",
2538=>x"00004",
2539=>x"00004",
2540=>x"00004",
2541=>x"00004",
2542=>x"00004",
2543=>x"00004",
2544=>x"00004",
2545=>x"00004",
2546=>x"00004",
2547=>x"00004",
2548=>x"00004",
2549=>x"00004",
2550=>x"00004",
2551=>x"00004",
2552=>x"00004",
2553=>x"00004",
2554=>x"00004",
2555=>x"00004",
2556=>x"00004",
2557=>x"00004",
2558=>x"00004",
2559=>x"00004",
2560=>x"00004",
2561=>x"00004",
2562=>x"00004",
2563=>x"00004",
2564=>x"00004",
2565=>x"00004",
2566=>x"00004",
2567=>x"00004",
2568=>x"00004",
2569=>x"00004",
2570=>x"00004",
2571=>x"00004",
2572=>x"00004",
2573=>x"00004",
2574=>x"00004",
2575=>x"00004",
2576=>x"00004",
2577=>x"00004",
2578=>x"00004",
2579=>x"00004",
2580=>x"00004",
2581=>x"00004",
2582=>x"00004",
2583=>x"00004",
2584=>x"00004",
2585=>x"00004",
2586=>x"00004",
2587=>x"00004",
2588=>x"00004",
2589=>x"00004",
2590=>x"00004",
2591=>x"00004",
2592=>x"00004",
2593=>x"00004",
2594=>x"00004",
2595=>x"00004",
2596=>x"00004",
2597=>x"00004",
2598=>x"00004",
2599=>x"00004",
2600=>x"00004",
2601=>x"00004",
2602=>x"00004",
2603=>x"00004",
2604=>x"00004",
2605=>x"00004",
2606=>x"00004",
2607=>x"00004",
2608=>x"00004",
2609=>x"00004",
2610=>x"00004",
2611=>x"00004",
2612=>x"00004",
2613=>x"00004",
2614=>x"00004",
2615=>x"00004",
2616=>x"00004",
2617=>x"00004",
2618=>x"00004",
2619=>x"00004",
2620=>x"00004",
2621=>x"00004",
2622=>x"00004",
2623=>x"00004",
2624=>x"00004",
2625=>x"00004",
2626=>x"00004",
2627=>x"00004",
2628=>x"00004",
2629=>x"00004",
2630=>x"00004",
2631=>x"00004",
2632=>x"00004",
2633=>x"00004",
2634=>x"00004",
2635=>x"00004",
2636=>x"00004",
2637=>x"00004",
2638=>x"00004",
2639=>x"00004",
2640=>x"00004",
2641=>x"00004",
2642=>x"00004",
2643=>x"00004",
2644=>x"00004",
2645=>x"00004",
2646=>x"00004",
2647=>x"00004",
2648=>x"00004",
2649=>x"00004",
2650=>x"00004",
2651=>x"00004",
2652=>x"00004",
2653=>x"00004",
2654=>x"00004",
2655=>x"00004",
2656=>x"00004",
2657=>x"00004",
2658=>x"00004",
2659=>x"00004",
2660=>x"00004",
2661=>x"00004",
2662=>x"00004",
2663=>x"00004",
2664=>x"00004",
2665=>x"00004",
2666=>x"00004",
2667=>x"00004",
2668=>x"00004",
2669=>x"00004",
2670=>x"00004",
2671=>x"00004",
2672=>x"00004",
2673=>x"00004",
2674=>x"00004",
2675=>x"00004",
2676=>x"00004",
2677=>x"00004",
2678=>x"00004",
2679=>x"00004",
2680=>x"00004",
2681=>x"00004",
2682=>x"00004",
2683=>x"00004",
2684=>x"00004",
2685=>x"00004",
2686=>x"00004",
2687=>x"00004",
2688=>x"00004",
2689=>x"00004",
2690=>x"00004",
2691=>x"00004",
2692=>x"00004",
2693=>x"00004",
2694=>x"00004",
2695=>x"00004",
2696=>x"00004",
2697=>x"00004",
2698=>x"00004",
2699=>x"00004",
2700=>x"00004",
2701=>x"00004",
2702=>x"00004",
2703=>x"00004",
2704=>x"00004",
2705=>x"00004",
2706=>x"00004",
2707=>x"00004",
2708=>x"00004",
2709=>x"00004",
2710=>x"00004",
2711=>x"00004",
2712=>x"00004",
2713=>x"00004",
2714=>x"00004",
2715=>x"00004",
2716=>x"00004",
2717=>x"00004",
2718=>x"00004",
2719=>x"00004",
2720=>x"00004",
2721=>x"00004",
2722=>x"00004",
2723=>x"00004",
2724=>x"00004",
2725=>x"00004",
2726=>x"00004",
2727=>x"00004",
2728=>x"00004",
2729=>x"00004",
2730=>x"00004",
2731=>x"00004",
2732=>x"00004",
2733=>x"00004",
2734=>x"00004",
2735=>x"00004",
2736=>x"00004",
2737=>x"00004",
2738=>x"00004",
2739=>x"00004",
2740=>x"00004",
2741=>x"00004",
2742=>x"00004",
2743=>x"00004",
2744=>x"00004",
2745=>x"00004",
2746=>x"00004",
2747=>x"00004",
2748=>x"00004",
2749=>x"00004",
2750=>x"00004",
2751=>x"00004",
2752=>x"00004",
2753=>x"00004",
2754=>x"00004",
2755=>x"00004",
2756=>x"00004",
2757=>x"00004",
2758=>x"00004",
2759=>x"00004",
2760=>x"00004",
2761=>x"00004",
2762=>x"00004",
2763=>x"00004",
2764=>x"00004",
2765=>x"00004",
2766=>x"00004",
2767=>x"00004",
2768=>x"00004",
2769=>x"00004",
2770=>x"00004",
2771=>x"00004",
2772=>x"00004",
2773=>x"00004",
2774=>x"00004",
2775=>x"00004",
2776=>x"00004",
2777=>x"00004",
2778=>x"00004",
2779=>x"00004",
2780=>x"00004",
2781=>x"00004",
2782=>x"00004",
2783=>x"00004",
2784=>x"00004",
2785=>x"00004",
2786=>x"00004",
2787=>x"00004",
2788=>x"00004",
2789=>x"00004",
2790=>x"00004",
2791=>x"00004",
2792=>x"00004",
2793=>x"00004",
2794=>x"00004",
2795=>x"00004",
2796=>x"00004",
2797=>x"00004",
2798=>x"00004",
2799=>x"00004",
2800=>x"00004",
2801=>x"00004",
2802=>x"00004",
2803=>x"00004",
2804=>x"00004",
2805=>x"00004",
2806=>x"00004",
2807=>x"00004",
2808=>x"00004",
2809=>x"00004",
2810=>x"00004",
2811=>x"00004",
2812=>x"00004",
2813=>x"00004",
2814=>x"00004",
2815=>x"00004",
2816=>x"00004",
2817=>x"00004",
2818=>x"00004",
2819=>x"00004",
2820=>x"00004",
2821=>x"00004",
2822=>x"00004",
2823=>x"00004",
2824=>x"00004",
2825=>x"00004",
2826=>x"00004",
2827=>x"00004",
2828=>x"00004",
2829=>x"00004",
2830=>x"00004",
2831=>x"00004",
2832=>x"00004",
2833=>x"00004",
2834=>x"00004",
2835=>x"00004",
2836=>x"00004",
2837=>x"00004",
2838=>x"00004",
2839=>x"00004",
2840=>x"00004",
2841=>x"00004",
2842=>x"00004",
2843=>x"00004",
2844=>x"00004",
2845=>x"00004",
2846=>x"00004",
2847=>x"00004",
2848=>x"00004",
2849=>x"00004",
2850=>x"00004",
2851=>x"00004",
2852=>x"00004",
2853=>x"00004",
2854=>x"00004",
2855=>x"00004",
2856=>x"00004",
2857=>x"00004",
2858=>x"00004",
2859=>x"00004",
2860=>x"00004",
2861=>x"00004",
2862=>x"00004",
2863=>x"00004",
2864=>x"00004",
2865=>x"00004",
2866=>x"00004",
2867=>x"00004",
2868=>x"00004",
2869=>x"00004",
2870=>x"00004",
2871=>x"00004",
2872=>x"00004",
2873=>x"00004",
2874=>x"00004",
2875=>x"00004",
2876=>x"00004",
2877=>x"00004",
2878=>x"00004",
2879=>x"00004",
2880=>x"00004",
2881=>x"00004",
2882=>x"00004",
2883=>x"00004",
2884=>x"00004",
2885=>x"00004",
2886=>x"00004",
2887=>x"00004",
2888=>x"00004",
2889=>x"00004",
2890=>x"00004",
2891=>x"00004",
2892=>x"00004",
2893=>x"00004",
2894=>x"00004",
2895=>x"00004",
2896=>x"00004",
2897=>x"00004",
2898=>x"00004",
2899=>x"00004",
2900=>x"00004",
2901=>x"00004",
2902=>x"00004",
2903=>x"00004",
2904=>x"00004",
2905=>x"00004",
2906=>x"00004",
2907=>x"00004",
2908=>x"00004",
2909=>x"00004",
2910=>x"00004",
2911=>x"00004",
2912=>x"00004",
2913=>x"00004",
2914=>x"00004",
2915=>x"00004",
2916=>x"00004",
2917=>x"00004",
2918=>x"00004",
2919=>x"00004",
2920=>x"00004",
2921=>x"00004",
2922=>x"00004",
2923=>x"00004",
2924=>x"00004",
2925=>x"00004",
2926=>x"00004",
2927=>x"00004",
2928=>x"00004",
2929=>x"00004",
2930=>x"00004",
2931=>x"00004",
2932=>x"00004",
2933=>x"00004",
2934=>x"00004",
2935=>x"00004",
2936=>x"00004",
2937=>x"00004",
2938=>x"00004",
2939=>x"00004",
2940=>x"00004",
2941=>x"00004",
2942=>x"00004",
2943=>x"00004",
2944=>x"00004",
2945=>x"00004",
2946=>x"00004",
2947=>x"00004",
2948=>x"00004",
2949=>x"00004",
2950=>x"00004",
2951=>x"00004",
2952=>x"00004",
2953=>x"00004",
2954=>x"00004",
2955=>x"00004",
2956=>x"00004",
2957=>x"00004",
2958=>x"00004",
2959=>x"00004",
2960=>x"00004",
2961=>x"00004",
2962=>x"00004",
2963=>x"00004",
2964=>x"00004",
2965=>x"00004",
2966=>x"00004",
2967=>x"00004",
2968=>x"00004",
2969=>x"00004",
2970=>x"00004",
2971=>x"00004",
2972=>x"00004",
2973=>x"00004",
2974=>x"00004",
2975=>x"00004",
2976=>x"00004",
2977=>x"00004",
2978=>x"00004",
2979=>x"00004",
2980=>x"00004",
2981=>x"00004",
2982=>x"00004",
2983=>x"00004",
2984=>x"00004",
2985=>x"00004",
2986=>x"00004",
2987=>x"00004",
2988=>x"00004",
2989=>x"00004",
2990=>x"00004",
2991=>x"00004",
2992=>x"00004",
2993=>x"00004",
2994=>x"00004",
2995=>x"00004",
2996=>x"00004",
2997=>x"00004",
2998=>x"00004",
2999=>x"00004",
3000=>x"00004",
3001=>x"00004",
3002=>x"00004",
3003=>x"00004",
3004=>x"00004",
3005=>x"00004",
3006=>x"00004",
3007=>x"00004",
3008=>x"00004",
3009=>x"00004",
3010=>x"00004",
3011=>x"00004",
3012=>x"00004",
3013=>x"00004",
3014=>x"00004",
3015=>x"00004",
3016=>x"00004",
3017=>x"00004",
3018=>x"00004",
3019=>x"00004",
3020=>x"00004",
3021=>x"00004",
3022=>x"00004",
3023=>x"00004",
3024=>x"00004",
3025=>x"00004",
3026=>x"00004",
3027=>x"00004",
3028=>x"00004",
3029=>x"00004",
3030=>x"00004",
3031=>x"00004",
3032=>x"00004",
3033=>x"00004",
3034=>x"00004",
3035=>x"00004",
3036=>x"00004",
3037=>x"00004",
3038=>x"00004",
3039=>x"00004",
3040=>x"00004",
3041=>x"00004",
3042=>x"00004",
3043=>x"00004",
3044=>x"00004",
3045=>x"00004",
3046=>x"00004",
3047=>x"00004",
3048=>x"00004",
3049=>x"00004",
3050=>x"00004",
3051=>x"00004",
3052=>x"00004",
3053=>x"00004",
3054=>x"00004",
3055=>x"00004",
3056=>x"00004",
3057=>x"00004",
3058=>x"00004",
3059=>x"00004",
3060=>x"00004",
3061=>x"00004",
3062=>x"00004",
3063=>x"00004",
3064=>x"00004",
3065=>x"00004",
3066=>x"00004",
3067=>x"00004",
3068=>x"00004",
3069=>x"00004",
3070=>x"00004",
3071=>x"00004",
3072=>x"00004",
3073=>x"00003",
3074=>x"00003",
3075=>x"00003",
3076=>x"00003",
3077=>x"00003",
3078=>x"00003",
3079=>x"00003",
3080=>x"00003",
3081=>x"00003",
3082=>x"00003",
3083=>x"00003",
3084=>x"00003",
3085=>x"00003",
3086=>x"00003",
3087=>x"00003",
3088=>x"00003",
3089=>x"00003",
3090=>x"00003",
3091=>x"00003",
3092=>x"00003",
3093=>x"00003",
3094=>x"00003",
3095=>x"00003",
3096=>x"00003",
3097=>x"00003",
3098=>x"00003",
3099=>x"00003",
3100=>x"00003",
3101=>x"00003",
3102=>x"00003",
3103=>x"00003",
3104=>x"00003",
3105=>x"00003",
3106=>x"00003",
3107=>x"00003",
3108=>x"00003",
3109=>x"00003",
3110=>x"00003",
3111=>x"00003",
3112=>x"00003",
3113=>x"00003",
3114=>x"00003",
3115=>x"00003",
3116=>x"00003",
3117=>x"00003",
3118=>x"00003",
3119=>x"00003",
3120=>x"00003",
3121=>x"00003",
3122=>x"00003",
3123=>x"00003",
3124=>x"00003",
3125=>x"00003",
3126=>x"00003",
3127=>x"00003",
3128=>x"00003",
3129=>x"00003",
3130=>x"00003",
3131=>x"00003",
3132=>x"00003",
3133=>x"00003",
3134=>x"00003",
3135=>x"00003",
3136=>x"00003",
3137=>x"00003",
3138=>x"00003",
3139=>x"00003",
3140=>x"00003",
3141=>x"00003",
3142=>x"00003",
3143=>x"00003",
3144=>x"00003",
3145=>x"00003",
3146=>x"00003",
3147=>x"00003",
3148=>x"00003",
3149=>x"00003",
3150=>x"00003",
3151=>x"00003",
3152=>x"00003",
3153=>x"00003",
3154=>x"00003",
3155=>x"00003",
3156=>x"00003",
3157=>x"00003",
3158=>x"00003",
3159=>x"00003",
3160=>x"00003",
3161=>x"00003",
3162=>x"00003",
3163=>x"00003",
3164=>x"00003",
3165=>x"00003",
3166=>x"00003",
3167=>x"00003",
3168=>x"00003",
3169=>x"00003",
3170=>x"00003",
3171=>x"00003",
3172=>x"00003",
3173=>x"00003",
3174=>x"00003",
3175=>x"00003",
3176=>x"00003",
3177=>x"00003",
3178=>x"00003",
3179=>x"00003",
3180=>x"00003",
3181=>x"00003",
3182=>x"00003",
3183=>x"00003",
3184=>x"00003",
3185=>x"00003",
3186=>x"00003",
3187=>x"00003",
3188=>x"00003",
3189=>x"00003",
3190=>x"00003",
3191=>x"00003",
3192=>x"00003",
3193=>x"00003",
3194=>x"00003",
3195=>x"00003",
3196=>x"00003",
3197=>x"00003",
3198=>x"00003",
3199=>x"00003",
3200=>x"00003",
3201=>x"00003",
3202=>x"00003",
3203=>x"00003",
3204=>x"00003",
3205=>x"00003",
3206=>x"00003",
3207=>x"00003",
3208=>x"00003",
3209=>x"00003",
3210=>x"00003",
3211=>x"00003",
3212=>x"00003",
3213=>x"00003",
3214=>x"00003",
3215=>x"00003",
3216=>x"00003",
3217=>x"00003",
3218=>x"00003",
3219=>x"00003",
3220=>x"00003",
3221=>x"00003",
3222=>x"00003",
3223=>x"00003",
3224=>x"00003",
3225=>x"00003",
3226=>x"00003",
3227=>x"00003",
3228=>x"00003",
3229=>x"00003",
3230=>x"00003",
3231=>x"00003",
3232=>x"00003",
3233=>x"00003",
3234=>x"00003",
3235=>x"00003",
3236=>x"00003",
3237=>x"00003",
3238=>x"00003",
3239=>x"00003",
3240=>x"00003",
3241=>x"00003",
3242=>x"00003",
3243=>x"00003",
3244=>x"00003",
3245=>x"00003",
3246=>x"00003",
3247=>x"00003",
3248=>x"00003",
3249=>x"00003",
3250=>x"00003",
3251=>x"00003",
3252=>x"00003",
3253=>x"00003",
3254=>x"00003",
3255=>x"00003",
3256=>x"00003",
3257=>x"00003",
3258=>x"00003",
3259=>x"00003",
3260=>x"00003",
3261=>x"00003",
3262=>x"00003",
3263=>x"00003",
3264=>x"00003",
3265=>x"00003",
3266=>x"00003",
3267=>x"00003",
3268=>x"00003",
3269=>x"00003",
3270=>x"00003",
3271=>x"00003",
3272=>x"00003",
3273=>x"00003",
3274=>x"00003",
3275=>x"00003",
3276=>x"00003",
3277=>x"00003",
3278=>x"00003",
3279=>x"00003",
3280=>x"00003",
3281=>x"00003",
3282=>x"00003",
3283=>x"00003",
3284=>x"00003",
3285=>x"00003",
3286=>x"00003",
3287=>x"00003",
3288=>x"00003",
3289=>x"00003",
3290=>x"00003",
3291=>x"00003",
3292=>x"00003",
3293=>x"00003",
3294=>x"00003",
3295=>x"00003",
3296=>x"00003",
3297=>x"00003",
3298=>x"00003",
3299=>x"00003",
3300=>x"00003",
3301=>x"00003",
3302=>x"00003",
3303=>x"00003",
3304=>x"00003",
3305=>x"00003",
3306=>x"00003",
3307=>x"00003",
3308=>x"00003",
3309=>x"00003",
3310=>x"00003",
3311=>x"00003",
3312=>x"00003",
3313=>x"00003",
3314=>x"00003",
3315=>x"00003",
3316=>x"00003",
3317=>x"00003",
3318=>x"00003",
3319=>x"00003",
3320=>x"00003",
3321=>x"00003",
3322=>x"00003",
3323=>x"00003",
3324=>x"00003",
3325=>x"00003",
3326=>x"00003",
3327=>x"00003",
3328=>x"00003",
3329=>x"00003",
3330=>x"00003",
3331=>x"00003",
3332=>x"00003",
3333=>x"00003",
3334=>x"00003",
3335=>x"00003",
3336=>x"00003",
3337=>x"00003",
3338=>x"00003",
3339=>x"00003",
3340=>x"00003",
3341=>x"00003",
3342=>x"00003",
3343=>x"00003",
3344=>x"00003",
3345=>x"00003",
3346=>x"00003",
3347=>x"00003",
3348=>x"00003",
3349=>x"00003",
3350=>x"00003",
3351=>x"00003",
3352=>x"00003",
3353=>x"00003",
3354=>x"00003",
3355=>x"00003",
3356=>x"00003",
3357=>x"00003",
3358=>x"00003",
3359=>x"00003",
3360=>x"00003",
3361=>x"00003",
3362=>x"00003",
3363=>x"00003",
3364=>x"00003",
3365=>x"00003",
3366=>x"00003",
3367=>x"00003",
3368=>x"00003",
3369=>x"00003",
3370=>x"00003",
3371=>x"00003",
3372=>x"00003",
3373=>x"00003",
3374=>x"00003",
3375=>x"00003",
3376=>x"00003",
3377=>x"00003",
3378=>x"00003",
3379=>x"00003",
3380=>x"00003",
3381=>x"00003",
3382=>x"00003",
3383=>x"00003",
3384=>x"00003",
3385=>x"00003",
3386=>x"00003",
3387=>x"00003",
3388=>x"00003",
3389=>x"00003",
3390=>x"00003",
3391=>x"00003",
3392=>x"00003",
3393=>x"00003",
3394=>x"00003",
3395=>x"00003",
3396=>x"00003",
3397=>x"00003",
3398=>x"00003",
3399=>x"00003",
3400=>x"00003",
3401=>x"00003",
3402=>x"00003",
3403=>x"00003",
3404=>x"00003",
3405=>x"00003",
3406=>x"00003",
3407=>x"00003",
3408=>x"00003",
3409=>x"00003",
3410=>x"00003",
3411=>x"00003",
3412=>x"00003",
3413=>x"00003",
3414=>x"00003",
3415=>x"00003",
3416=>x"00003",
3417=>x"00003",
3418=>x"00003",
3419=>x"00003",
3420=>x"00003",
3421=>x"00003",
3422=>x"00003",
3423=>x"00003",
3424=>x"00003",
3425=>x"00003",
3426=>x"00003",
3427=>x"00003",
3428=>x"00003",
3429=>x"00003",
3430=>x"00003",
3431=>x"00003",
3432=>x"00003",
3433=>x"00003",
3434=>x"00003",
3435=>x"00003",
3436=>x"00003",
3437=>x"00003",
3438=>x"00003",
3439=>x"00003",
3440=>x"00003",
3441=>x"00003",
3442=>x"00003",
3443=>x"00003",
3444=>x"00003",
3445=>x"00003",
3446=>x"00003",
3447=>x"00003",
3448=>x"00003",
3449=>x"00003",
3450=>x"00003",
3451=>x"00003",
3452=>x"00003",
3453=>x"00003",
3454=>x"00003",
3455=>x"00003",
3456=>x"00003",
3457=>x"00003",
3458=>x"00003",
3459=>x"00003",
3460=>x"00003",
3461=>x"00003",
3462=>x"00003",
3463=>x"00003",
3464=>x"00003",
3465=>x"00003",
3466=>x"00003",
3467=>x"00003",
3468=>x"00003",
3469=>x"00003",
3470=>x"00003",
3471=>x"00003",
3472=>x"00003",
3473=>x"00003",
3474=>x"00003",
3475=>x"00003",
3476=>x"00003",
3477=>x"00003",
3478=>x"00003",
3479=>x"00003",
3480=>x"00003",
3481=>x"00003",
3482=>x"00003",
3483=>x"00003",
3484=>x"00003",
3485=>x"00003",
3486=>x"00003",
3487=>x"00003",
3488=>x"00003",
3489=>x"00003",
3490=>x"00003",
3491=>x"00003",
3492=>x"00003",
3493=>x"00003",
3494=>x"00003",
3495=>x"00003",
3496=>x"00003",
3497=>x"00003",
3498=>x"00003",
3499=>x"00003",
3500=>x"00003",
3501=>x"00003",
3502=>x"00003",
3503=>x"00003",
3504=>x"00003",
3505=>x"00003",
3506=>x"00003",
3507=>x"00003",
3508=>x"00003",
3509=>x"00003",
3510=>x"00003",
3511=>x"00003",
3512=>x"00003",
3513=>x"00003",
3514=>x"00003",
3515=>x"00003",
3516=>x"00003",
3517=>x"00003",
3518=>x"00003",
3519=>x"00003",
3520=>x"00003",
3521=>x"00003",
3522=>x"00003",
3523=>x"00003",
3524=>x"00003",
3525=>x"00003",
3526=>x"00003",
3527=>x"00003",
3528=>x"00003",
3529=>x"00003",
3530=>x"00003",
3531=>x"00003",
3532=>x"00003",
3533=>x"00003",
3534=>x"00003",
3535=>x"00003",
3536=>x"00003",
3537=>x"00003",
3538=>x"00003",
3539=>x"00003",
3540=>x"00003",
3541=>x"00003",
3542=>x"00003",
3543=>x"00003",
3544=>x"00003",
3545=>x"00003",
3546=>x"00003",
3547=>x"00003",
3548=>x"00003",
3549=>x"00003",
3550=>x"00003",
3551=>x"00003",
3552=>x"00003",
3553=>x"00003",
3554=>x"00003",
3555=>x"00003",
3556=>x"00003",
3557=>x"00003",
3558=>x"00003",
3559=>x"00003",
3560=>x"00003",
3561=>x"00003",
3562=>x"00003",
3563=>x"00003",
3564=>x"00003",
3565=>x"00003",
3566=>x"00003",
3567=>x"00003",
3568=>x"00003",
3569=>x"00003",
3570=>x"00003",
3571=>x"00003",
3572=>x"00003",
3573=>x"00003",
3574=>x"00003",
3575=>x"00003",
3576=>x"00003",
3577=>x"00003",
3578=>x"00003",
3579=>x"00003",
3580=>x"00003",
3581=>x"00003",
3582=>x"00003",
3583=>x"00003",
3584=>x"00003",
3585=>x"00003",
3586=>x"00003",
3587=>x"00003",
3588=>x"00003",
3589=>x"00003",
3590=>x"00003",
3591=>x"00003",
3592=>x"00003",
3593=>x"00003",
3594=>x"00003",
3595=>x"00003",
3596=>x"00003",
3597=>x"00003",
3598=>x"00003",
3599=>x"00003",
3600=>x"00003",
3601=>x"00003",
3602=>x"00003",
3603=>x"00003",
3604=>x"00003",
3605=>x"00003",
3606=>x"00003",
3607=>x"00003",
3608=>x"00003",
3609=>x"00003",
3610=>x"00003",
3611=>x"00003",
3612=>x"00003",
3613=>x"00003",
3614=>x"00003",
3615=>x"00003",
3616=>x"00003",
3617=>x"00003",
3618=>x"00003",
3619=>x"00003",
3620=>x"00003",
3621=>x"00003",
3622=>x"00003",
3623=>x"00003",
3624=>x"00003",
3625=>x"00003",
3626=>x"00003",
3627=>x"00003",
3628=>x"00003",
3629=>x"00003",
3630=>x"00003",
3631=>x"00003",
3632=>x"00003",
3633=>x"00003",
3634=>x"00003",
3635=>x"00003",
3636=>x"00003",
3637=>x"00003",
3638=>x"00003",
3639=>x"00003",
3640=>x"00003",
3641=>x"00003",
3642=>x"00003",
3643=>x"00003",
3644=>x"00003",
3645=>x"00003",
3646=>x"00003",
3647=>x"00003",
3648=>x"00003",
3649=>x"00003",
3650=>x"00003",
3651=>x"00003",
3652=>x"00003",
3653=>x"00003",
3654=>x"00003",
3655=>x"00003",
3656=>x"00003",
3657=>x"00003",
3658=>x"00003",
3659=>x"00003",
3660=>x"00003",
3661=>x"00003",
3662=>x"00003",
3663=>x"00003",
3664=>x"00003",
3665=>x"00003",
3666=>x"00003",
3667=>x"00003",
3668=>x"00003",
3669=>x"00003",
3670=>x"00003",
3671=>x"00003",
3672=>x"00003",
3673=>x"00003",
3674=>x"00003",
3675=>x"00003",
3676=>x"00003",
3677=>x"00003",
3678=>x"00003",
3679=>x"00003",
3680=>x"00003",
3681=>x"00003",
3682=>x"00003",
3683=>x"00003",
3684=>x"00003",
3685=>x"00003",
3686=>x"00003",
3687=>x"00003",
3688=>x"00003",
3689=>x"00003",
3690=>x"00003",
3691=>x"00003",
3692=>x"00003",
3693=>x"00003",
3694=>x"00003",
3695=>x"00003",
3696=>x"00003",
3697=>x"00003",
3698=>x"00003",
3699=>x"00003",
3700=>x"00003",
3701=>x"00003",
3702=>x"00003",
3703=>x"00003",
3704=>x"00003",
3705=>x"00003",
3706=>x"00003",
3707=>x"00003",
3708=>x"00003",
3709=>x"00003",
3710=>x"00003",
3711=>x"00003",
3712=>x"00003",
3713=>x"00003",
3714=>x"00003",
3715=>x"00003",
3716=>x"00003",
3717=>x"00003",
3718=>x"00003",
3719=>x"00003",
3720=>x"00003",
3721=>x"00003",
3722=>x"00003",
3723=>x"00003",
3724=>x"00003",
3725=>x"00003",
3726=>x"00003",
3727=>x"00003",
3728=>x"00003",
3729=>x"00003",
3730=>x"00003",
3731=>x"00003",
3732=>x"00003",
3733=>x"00003",
3734=>x"00003",
3735=>x"00003",
3736=>x"00003",
3737=>x"00003",
3738=>x"00003",
3739=>x"00003",
3740=>x"00003",
3741=>x"00003",
3742=>x"00003",
3743=>x"00003",
3744=>x"00003",
3745=>x"00003",
3746=>x"00003",
3747=>x"00003",
3748=>x"00003",
3749=>x"00003",
3750=>x"00003",
3751=>x"00003",
3752=>x"00003",
3753=>x"00003",
3754=>x"00003",
3755=>x"00003",
3756=>x"00003",
3757=>x"00003",
3758=>x"00003",
3759=>x"00003",
3760=>x"00003",
3761=>x"00003",
3762=>x"00003",
3763=>x"00003",
3764=>x"00003",
3765=>x"00003",
3766=>x"00003",
3767=>x"00003",
3768=>x"00003",
3769=>x"00003",
3770=>x"00003",
3771=>x"00003",
3772=>x"00003",
3773=>x"00003",
3774=>x"00003",
3775=>x"00003",
3776=>x"00003",
3777=>x"00003",
3778=>x"00003",
3779=>x"00003",
3780=>x"00003",
3781=>x"00003",
3782=>x"00003",
3783=>x"00003",
3784=>x"00003",
3785=>x"00003",
3786=>x"00003",
3787=>x"00003",
3788=>x"00003",
3789=>x"00003",
3790=>x"00003",
3791=>x"00003",
3792=>x"00003",
3793=>x"00003",
3794=>x"00003",
3795=>x"00003",
3796=>x"00003",
3797=>x"00003",
3798=>x"00003",
3799=>x"00003",
3800=>x"00003",
3801=>x"00003",
3802=>x"00003",
3803=>x"00003",
3804=>x"00003",
3805=>x"00003",
3806=>x"00003",
3807=>x"00003",
3808=>x"00003",
3809=>x"00003",
3810=>x"00003",
3811=>x"00003",
3812=>x"00003",
3813=>x"00003",
3814=>x"00003",
3815=>x"00003",
3816=>x"00003",
3817=>x"00003",
3818=>x"00003",
3819=>x"00003",
3820=>x"00003",
3821=>x"00003",
3822=>x"00003",
3823=>x"00003",
3824=>x"00003",
3825=>x"00003",
3826=>x"00003",
3827=>x"00003",
3828=>x"00003",
3829=>x"00003",
3830=>x"00003",
3831=>x"00003",
3832=>x"00003",
3833=>x"00003",
3834=>x"00003",
3835=>x"00003",
3836=>x"00003",
3837=>x"00003",
3838=>x"00003",
3839=>x"00003",
3840=>x"00003",
3841=>x"00003",
3842=>x"00003",
3843=>x"00003",
3844=>x"00003",
3845=>x"00003",
3846=>x"00003",
3847=>x"00003",
3848=>x"00003",
3849=>x"00003",
3850=>x"00003",
3851=>x"00003",
3852=>x"00003",
3853=>x"00003",
3854=>x"00003",
3855=>x"00003",
3856=>x"00003",
3857=>x"00003",
3858=>x"00003",
3859=>x"00003",
3860=>x"00003",
3861=>x"00003",
3862=>x"00003",
3863=>x"00003",
3864=>x"00003",
3865=>x"00003",
3866=>x"00003",
3867=>x"00003",
3868=>x"00003",
3869=>x"00003",
3870=>x"00003",
3871=>x"00003",
3872=>x"00003",
3873=>x"00003",
3874=>x"00003",
3875=>x"00003",
3876=>x"00003",
3877=>x"00003",
3878=>x"00003",
3879=>x"00003",
3880=>x"00003",
3881=>x"00003",
3882=>x"00003",
3883=>x"00003",
3884=>x"00003",
3885=>x"00003",
3886=>x"00003",
3887=>x"00003",
3888=>x"00003",
3889=>x"00003",
3890=>x"00003",
3891=>x"00003",
3892=>x"00003",
3893=>x"00003",
3894=>x"00003",
3895=>x"00003",
3896=>x"00003",
3897=>x"00003",
3898=>x"00003",
3899=>x"00003",
3900=>x"00003",
3901=>x"00003",
3902=>x"00003",
3903=>x"00003",
3904=>x"00003",
3905=>x"00003",
3906=>x"00003",
3907=>x"00003",
3908=>x"00003",
3909=>x"00003",
3910=>x"00003",
3911=>x"00003",
3912=>x"00003",
3913=>x"00003",
3914=>x"00003",
3915=>x"00003",
3916=>x"00003",
3917=>x"00003",
3918=>x"00003",
3919=>x"00003",
3920=>x"00003",
3921=>x"00003",
3922=>x"00003",
3923=>x"00003",
3924=>x"00003",
3925=>x"00003",
3926=>x"00003",
3927=>x"00003",
3928=>x"00003",
3929=>x"00003",
3930=>x"00003",
3931=>x"00003",
3932=>x"00003",
3933=>x"00003",
3934=>x"00003",
3935=>x"00003",
3936=>x"00003",
3937=>x"00003",
3938=>x"00003",
3939=>x"00003",
3940=>x"00003",
3941=>x"00003",
3942=>x"00003",
3943=>x"00003",
3944=>x"00003",
3945=>x"00003",
3946=>x"00003",
3947=>x"00003",
3948=>x"00003",
3949=>x"00003",
3950=>x"00003",
3951=>x"00003",
3952=>x"00003",
3953=>x"00003",
3954=>x"00003",
3955=>x"00003",
3956=>x"00003",
3957=>x"00003",
3958=>x"00003",
3959=>x"00003",
3960=>x"00003",
3961=>x"00003",
3962=>x"00003",
3963=>x"00003",
3964=>x"00003",
3965=>x"00003",
3966=>x"00003",
3967=>x"00003",
3968=>x"00003",
3969=>x"00003",
3970=>x"00003",
3971=>x"00003",
3972=>x"00003",
3973=>x"00003",
3974=>x"00003",
3975=>x"00003",
3976=>x"00003",
3977=>x"00003",
3978=>x"00003",
3979=>x"00003",
3980=>x"00003",
3981=>x"00003",
3982=>x"00003",
3983=>x"00003",
3984=>x"00003",
3985=>x"00003",
3986=>x"00003",
3987=>x"00003",
3988=>x"00003",
3989=>x"00003",
3990=>x"00003",
3991=>x"00003",
3992=>x"00003",
3993=>x"00003",
3994=>x"00003",
3995=>x"00003",
3996=>x"00003",
3997=>x"00003",
3998=>x"00003",
3999=>x"00003",
4000=>x"00003",
4001=>x"00003",
4002=>x"00003",
4003=>x"00003",
4004=>x"00003",
4005=>x"00003",
4006=>x"00003",
4007=>x"00003",
4008=>x"00003",
4009=>x"00003",
4010=>x"00003",
4011=>x"00003",
4012=>x"00003",
4013=>x"00003",
4014=>x"00003",
4015=>x"00003",
4016=>x"00003",
4017=>x"00003",
4018=>x"00003",
4019=>x"00003",
4020=>x"00003",
4021=>x"00003",
4022=>x"00003",
4023=>x"00003",
4024=>x"00003",
4025=>x"00003",
4026=>x"00003",
4027=>x"00003",
4028=>x"00003",
4029=>x"00003",
4030=>x"00003",
4031=>x"00003",
4032=>x"00003",
4033=>x"00003",
4034=>x"00003",
4035=>x"00003",
4036=>x"00003",
4037=>x"00003",
4038=>x"00003",
4039=>x"00003",
4040=>x"00003",
4041=>x"00003",
4042=>x"00003",
4043=>x"00003",
4044=>x"00003",
4045=>x"00003",
4046=>x"00003",
4047=>x"00003",
4048=>x"00003",
4049=>x"00003",
4050=>x"00003",
4051=>x"00003",
4052=>x"00003",
4053=>x"00003",
4054=>x"00003",
4055=>x"00003",
4056=>x"00003",
4057=>x"00003",
4058=>x"00003",
4059=>x"00003",
4060=>x"00003",
4061=>x"00003",
4062=>x"00003",
4063=>x"00003",
4064=>x"00003",
4065=>x"00003",
4066=>x"00003",
4067=>x"00003",
4068=>x"00003",
4069=>x"00003",
4070=>x"00003",
4071=>x"00003",
4072=>x"00003",
4073=>x"00003",
4074=>x"00003",
4075=>x"00003",
4076=>x"00003",
4077=>x"00003",
4078=>x"00003",
4079=>x"00003",
4080=>x"00003",
4081=>x"00003",
4082=>x"00003",
4083=>x"00003",
4084=>x"00003",
4085=>x"00003",
4086=>x"00003",
4087=>x"00003",
4088=>x"00003",
4089=>x"00003",
4090=>x"00003",
4091=>x"00003",
4092=>x"00003",
4093=>x"00003",
4094=>x"00003",

others=>x"00000"
);
begin
Cout<=memory(to_integer(unsigned(addr)));

end Behavioral;