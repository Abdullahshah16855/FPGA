library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.ALL;

entity ROM_L is
    Port ( addr : in STD_LOGIC_VECTOR (39 downto 0);
           Cout : out STD_LOGIC_VECTOR (19 downto 0));
end ROM_L;

architecture Behavioral of ROM_L is
type vector is Array(0 to 15000) of Std_logic_vector(19 downto 0);
Constant memory: vector:=
(0=>x"00000",
1=>x"00000",
2=>x"00000",
3=>x"00000",
4=>x"00000",
5=>x"00000",
6=>x"00000",
7=>x"00000",
8=>x"00000",
9=>x"00000",
10=>x"00000",
11=>x"00000",
12=>x"00000",
13=>x"00000",
14=>x"00001",
15=>x"00001",
16=>x"00001",
17=>x"00001",
18=>x"00001",
19=>x"00001",
20=>x"00001",
21=>x"00001",
22=>x"00001",
23=>x"00001",
24=>x"00001",
25=>x"00001",
26=>x"00001",
27=>x"00001",
28=>x"00002",
29=>x"00002",
30=>x"00002",
31=>x"00002",
32=>x"00002",
33=>x"00002",
34=>x"00002",
35=>x"00002",
36=>x"00002",
37=>x"00002",
38=>x"00002",
39=>x"00002",
40=>x"00002",
41=>x"00002",
42=>x"00003",
43=>x"00003",
44=>x"00003",
45=>x"00003",
46=>x"00003",
47=>x"00003",
48=>x"00003",
49=>x"00003",
50=>x"00003",
51=>x"00003",
52=>x"00003",
53=>x"00003",
54=>x"00003",
55=>x"00003",
56=>x"00004",
57=>x"00004",
58=>x"00004",
59=>x"00004",
60=>x"00004",
61=>x"00004",
62=>x"00004",
63=>x"00004",
64=>x"00004",
65=>x"00004",
66=>x"00004",
67=>x"00004",
68=>x"00004",
69=>x"00004",
70=>x"00005",
71=>x"00005",
72=>x"00005",
73=>x"00005",
74=>x"00005",
75=>x"00005",
76=>x"00005",
77=>x"00005",
78=>x"00005",
79=>x"00005",
80=>x"00005",
81=>x"00005",
82=>x"00005",
83=>x"00005",
84=>x"00006",
85=>x"00006",
86=>x"00006",
87=>x"00006",
88=>x"00006",
89=>x"00006",
90=>x"00006",
91=>x"00006",
92=>x"00006",
93=>x"00006",
94=>x"00006",
95=>x"00006",
96=>x"00006",
97=>x"00006",
98=>x"00007",
99=>x"00007",
100=>x"00007",
101=>x"00007",
102=>x"00007",
103=>x"00007",
104=>x"00007",
105=>x"00007",
106=>x"00007",
107=>x"00007",
108=>x"00007",
109=>x"00007",
110=>x"00007",
111=>x"00007",
112=>x"00008",
113=>x"00008",
114=>x"00008",
115=>x"00008",
116=>x"00008",
117=>x"00008",
118=>x"00008",
119=>x"00008",
120=>x"00008",
121=>x"00008",
122=>x"00008",
123=>x"00008",
124=>x"00008",
125=>x"00008",
126=>x"00009",
127=>x"00009",
128=>x"00009",
129=>x"00009",
130=>x"00009",
131=>x"00009",
132=>x"00009",
133=>x"00009",
134=>x"00009",
135=>x"00009",
136=>x"00009",
137=>x"00009",
138=>x"00009",
139=>x"00009",
140=>x"0000a",
141=>x"0000a",
142=>x"0000a",
143=>x"0000a",
144=>x"0000a",
145=>x"0000a",
146=>x"0000a",
147=>x"0000a",
148=>x"0000a",
149=>x"0000a",
150=>x"0000a",
151=>x"0000a",
152=>x"0000a",
153=>x"0000a",
154=>x"0000b",
155=>x"0000b",
156=>x"0000b",
157=>x"0000b",
158=>x"0000b",
159=>x"0000b",
160=>x"0000b",
161=>x"0000b",
162=>x"0000b",
163=>x"0000b",
164=>x"0000b",
165=>x"0000b",
166=>x"0000b",
167=>x"0000b",
168=>x"0000c",
169=>x"0000c",
170=>x"0000c",
171=>x"0000c",
172=>x"0000c",
173=>x"0000c",
174=>x"0000c",
175=>x"0000c",
176=>x"0000c",
177=>x"0000c",
178=>x"0000c",
179=>x"0000c",
180=>x"0000c",
181=>x"0000c",
182=>x"0000d",
183=>x"0000d",
184=>x"0000d",
185=>x"0000d",
186=>x"0000d",
187=>x"0000d",
188=>x"0000d",
189=>x"0000d",
190=>x"0000d",
191=>x"0000d",
192=>x"0000d",
193=>x"0000d",
194=>x"0000d",
195=>x"0000d",
196=>x"0000e",
197=>x"0000e",
198=>x"0000e",
199=>x"0000e",
200=>x"0000e",
201=>x"0000e",
202=>x"0000e",
203=>x"0000e",
204=>x"0000e",
205=>x"0000e",
206=>x"0000e",
207=>x"0000e",
208=>x"0000e",
209=>x"0000e",
210=>x"0000f",
211=>x"0000f",
212=>x"0000f",
213=>x"0000f",
214=>x"0000f",
215=>x"0000f",
216=>x"0000f",
217=>x"0000f",
218=>x"0000f",
219=>x"0000f",
220=>x"0000f",
221=>x"0000f",
222=>x"0000f",
223=>x"0000f",
224=>x"00010",
225=>x"00010",
226=>x"00010",
227=>x"00010",
228=>x"00010",
229=>x"00010",
230=>x"00010",
231=>x"00010",
232=>x"00010",
233=>x"00010",
234=>x"00010",
235=>x"00010",
236=>x"00010",
237=>x"00010",
238=>x"00011",
239=>x"00011",
240=>x"00011",
241=>x"00011",
242=>x"00011",
243=>x"00011",
244=>x"00011",
245=>x"00011",
246=>x"00011",
247=>x"00011",
248=>x"00011",
249=>x"00011",
250=>x"00011",
251=>x"00011",
252=>x"00012",
253=>x"00012",
254=>x"00012",
255=>x"00012",
256=>x"00012",
257=>x"00012",
258=>x"00012",
259=>x"00012",
260=>x"00012",
261=>x"00012",
262=>x"00012",
263=>x"00012",
264=>x"00012",
265=>x"00012",
266=>x"00013",
267=>x"00013",
268=>x"00013",
269=>x"00013",
270=>x"00013",
271=>x"00013",
272=>x"00013",
273=>x"00013",
274=>x"00013",
275=>x"00013",
276=>x"00013",
277=>x"00013",
278=>x"00013",
279=>x"00013",
280=>x"00014",
281=>x"00014",
282=>x"00014",
283=>x"00014",
284=>x"00014",
285=>x"00014",
286=>x"00014",
287=>x"00014",
288=>x"00014",
289=>x"00014",
290=>x"00014",
291=>x"00014",
292=>x"00014",
293=>x"00014",
294=>x"00015",
295=>x"00015",
296=>x"00015",
297=>x"00015",
298=>x"00015",
299=>x"00015",
300=>x"00015",
301=>x"00015",
302=>x"00015",
303=>x"00015",
304=>x"00015",
305=>x"00015",
306=>x"00015",
307=>x"00015",
308=>x"00016",
309=>x"00016",
310=>x"00016",
311=>x"00016",
312=>x"00016",
313=>x"00016",
314=>x"00016",
315=>x"00016",
316=>x"00016",
317=>x"00016",
318=>x"00016",
319=>x"00016",
320=>x"00016",
321=>x"00016",
322=>x"00017",
323=>x"00017",
324=>x"00017",
325=>x"00017",
326=>x"00017",
327=>x"00017",
328=>x"00017",
329=>x"00017",
330=>x"00017",
331=>x"00017",
332=>x"00017",
333=>x"00017",
334=>x"00017",
335=>x"00017",
336=>x"00018",
337=>x"00018",
338=>x"00018",
339=>x"00018",
340=>x"00018",
341=>x"00018",
342=>x"00018",
343=>x"00018",
344=>x"00018",
345=>x"00018",
346=>x"00018",
347=>x"00018",
348=>x"00018",
349=>x"00018",
350=>x"00019",
351=>x"00019",
352=>x"00019",
353=>x"00019",
354=>x"00019",
355=>x"00019",
356=>x"00019",
357=>x"00019",
358=>x"00019",
359=>x"00019",
360=>x"00019",
361=>x"00019",
362=>x"00019",
363=>x"00019",
364=>x"0001a",
365=>x"0001a",
366=>x"0001a",
367=>x"0001a",
368=>x"0001a",
369=>x"0001a",
370=>x"0001a",
371=>x"0001a",
372=>x"0001a",
373=>x"0001a",
374=>x"0001a",
375=>x"0001a",
376=>x"0001a",
377=>x"0001a",
378=>x"0001b",
379=>x"0001b",
380=>x"0001b",
381=>x"0001b",
382=>x"0001b",
383=>x"0001b",
384=>x"0001b",
385=>x"0001b",
386=>x"0001b",
387=>x"0001b",
388=>x"0001b",
389=>x"0001b",
390=>x"0001b",
391=>x"0001b",
392=>x"0001c",
393=>x"0001c",
394=>x"0001c",
395=>x"0001c",
396=>x"0001c",
397=>x"0001c",
398=>x"0001c",
399=>x"0001c",
400=>x"0001c",
401=>x"0001c",
402=>x"0001c",
403=>x"0001c",
404=>x"0001c",
405=>x"0001c",
406=>x"0001d",
407=>x"0001d",
408=>x"0001d",
409=>x"0001d",
410=>x"0001d",
411=>x"0001d",
412=>x"0001d",
413=>x"0001d",
414=>x"0001d",
415=>x"0001d",
416=>x"0001d",
417=>x"0001d",
418=>x"0001d",
419=>x"0001d",
420=>x"0001e",
421=>x"0001e",
422=>x"0001e",
423=>x"0001e",
424=>x"0001e",
425=>x"0001e",
426=>x"0001e",
427=>x"0001e",
428=>x"0001e",
429=>x"0001e",
430=>x"0001e",
431=>x"0001e",
432=>x"0001e",
433=>x"0001e",
434=>x"0001f",
435=>x"0001f",
436=>x"0001f",
437=>x"0001f",
438=>x"0001f",
439=>x"0001f",
440=>x"0001f",
441=>x"0001f",
442=>x"0001f",
443=>x"0001f",
444=>x"0001f",
445=>x"0001f",
446=>x"0001f",
447=>x"0001f",
448=>x"00020",
449=>x"00020",
450=>x"00020",
451=>x"00020",
452=>x"00020",
453=>x"00020",
454=>x"00020",
455=>x"00020",
456=>x"00020",
457=>x"00020",
458=>x"00020",
459=>x"00020",
460=>x"00020",
461=>x"00020",
462=>x"00021",
463=>x"00021",
464=>x"00021",
465=>x"00021",
466=>x"00021",
467=>x"00021",
468=>x"00021",
469=>x"00021",
470=>x"00021",
471=>x"00021",
472=>x"00021",
473=>x"00021",
474=>x"00021",
475=>x"00021",
476=>x"00022",
477=>x"00022",
478=>x"00022",
479=>x"00022",
480=>x"00022",
481=>x"00022",
482=>x"00022",
483=>x"00022",
484=>x"00022",
485=>x"00022",
486=>x"00022",
487=>x"00022",
488=>x"00022",
489=>x"00022",
490=>x"00023",
491=>x"00023",
492=>x"00023",
493=>x"00023",
494=>x"00023",
495=>x"00023",
496=>x"00023",
497=>x"00023",
498=>x"00023",
499=>x"00023",
500=>x"00023",
501=>x"00023",
502=>x"00023",
503=>x"00023",
504=>x"00024",
505=>x"00024",
506=>x"00024",
507=>x"00024",
508=>x"00024",
509=>x"00024",
510=>x"00024",
511=>x"00024",
512=>x"00024",
513=>x"00024",
514=>x"00024",
515=>x"00024",
516=>x"00024",
517=>x"00024",
518=>x"00025",
519=>x"00025",
520=>x"00025",
521=>x"00025",
522=>x"00025",
523=>x"00025",
524=>x"00025",
525=>x"00025",
526=>x"00025",
527=>x"00025",
528=>x"00025",
529=>x"00025",
530=>x"00025",
531=>x"00025",
532=>x"00026",
533=>x"00026",
534=>x"00026",
535=>x"00026",
536=>x"00026",
537=>x"00026",
538=>x"00026",
539=>x"00026",
540=>x"00026",
541=>x"00026",
542=>x"00026",
543=>x"00026",
544=>x"00026",
545=>x"00026",
546=>x"00027",
547=>x"00027",
548=>x"00027",
549=>x"00027",
550=>x"00027",
551=>x"00027",
552=>x"00027",
553=>x"00027",
554=>x"00027",
555=>x"00027",
556=>x"00027",
557=>x"00027",
558=>x"00027",
559=>x"00027",
560=>x"00028",
561=>x"00028",
562=>x"00028",
563=>x"00028",
564=>x"00028",
565=>x"00028",
566=>x"00028",
567=>x"00028",
568=>x"00028",
569=>x"00028",
570=>x"00028",
571=>x"00028",
572=>x"00028",
573=>x"00028",
574=>x"00029",
575=>x"00029",
576=>x"00029",
577=>x"00029",
578=>x"00029",
579=>x"00029",
580=>x"00029",
581=>x"00029",
582=>x"00029",
583=>x"00029",
584=>x"00029",
585=>x"00029",
586=>x"00029",
587=>x"00029",
588=>x"0002a",
589=>x"0002a",
590=>x"0002a",
591=>x"0002a",
592=>x"0002a",
593=>x"0002a",
594=>x"0002a",
595=>x"0002a",
596=>x"0002a",
597=>x"0002a",
598=>x"0002a",
599=>x"0002a",
600=>x"0002a",
601=>x"0002a",
602=>x"0002b",
603=>x"0002b",
604=>x"0002b",
605=>x"0002b",
606=>x"0002b",
607=>x"0002b",
608=>x"0002b",
609=>x"0002b",
610=>x"0002b",
611=>x"0002b",
612=>x"0002b",
613=>x"0002b",
614=>x"0002b",
615=>x"0002b",
616=>x"0002c",
617=>x"0002c",
618=>x"0002c",
619=>x"0002c",
620=>x"0002c",
621=>x"0002c",
622=>x"0002c",
623=>x"0002c",
624=>x"0002c",
625=>x"0002c",
626=>x"0002c",
627=>x"0002c",
628=>x"0002c",
629=>x"0002c",
630=>x"0002d",
631=>x"0002d",
632=>x"0002d",
633=>x"0002d",
634=>x"0002d",
635=>x"0002d",
636=>x"0002d",
637=>x"0002d",
638=>x"0002d",
639=>x"0002d",
640=>x"0002d",
641=>x"0002d",
642=>x"0002d",
643=>x"0002d",
644=>x"0002e",
645=>x"0002e",
646=>x"0002e",
647=>x"0002e",
648=>x"0002e",
649=>x"0002e",
650=>x"0002e",
651=>x"0002e",
652=>x"0002e",
653=>x"0002e",
654=>x"0002e",
655=>x"0002e",
656=>x"0002e",
657=>x"0002e",
658=>x"0002f",
659=>x"0002f",
660=>x"0002f",
661=>x"0002f",
662=>x"0002f",
663=>x"0002f",
664=>x"0002f",
665=>x"0002f",
666=>x"0002f",
667=>x"0002f",
668=>x"0002f",
669=>x"0002f",
670=>x"0002f",
671=>x"0002f",
672=>x"00030",
673=>x"00030",
674=>x"00030",
675=>x"00030",
676=>x"00030",
677=>x"00030",
678=>x"00030",
679=>x"00030",
680=>x"00030",
681=>x"00030",
682=>x"00030",
683=>x"00030",
684=>x"00030",
685=>x"00030",
686=>x"00031",
687=>x"00031",
688=>x"00031",
689=>x"00031",
690=>x"00031",
691=>x"00031",
692=>x"00031",
693=>x"00031",
694=>x"00031",
695=>x"00031",
696=>x"00031",
697=>x"00031",
698=>x"00031",
699=>x"00031",
700=>x"00032",
701=>x"00032",
702=>x"00032",
703=>x"00032",
704=>x"00032",
705=>x"00032",
706=>x"00032",
707=>x"00032",
708=>x"00032",
709=>x"00032",
710=>x"00032",
711=>x"00032",
712=>x"00032",
713=>x"00032",
714=>x"00033",
715=>x"00033",
716=>x"00033",
717=>x"00033",
718=>x"00033",
719=>x"00033",
720=>x"00033",
721=>x"00033",
722=>x"00033",
723=>x"00033",
724=>x"00033",
725=>x"00033",
726=>x"00033",
727=>x"00033",
728=>x"00034",
729=>x"00034",
730=>x"00034",
731=>x"00034",
732=>x"00034",
733=>x"00034",
734=>x"00034",
735=>x"00034",
736=>x"00034",
737=>x"00034",
738=>x"00034",
739=>x"00034",
740=>x"00034",
741=>x"00034",
742=>x"00035",
743=>x"00035",
744=>x"00035",
745=>x"00035",
746=>x"00035",
747=>x"00035",
748=>x"00035",
749=>x"00035",
750=>x"00035",
751=>x"00035",
752=>x"00035",
753=>x"00035",
754=>x"00035",
755=>x"00035",
756=>x"00036",
757=>x"00036",
758=>x"00036",
759=>x"00036",
760=>x"00036",
761=>x"00036",
762=>x"00036",
763=>x"00036",
764=>x"00036",
765=>x"00036",
766=>x"00036",
767=>x"00036",
768=>x"00036",
769=>x"00036",
770=>x"00037",
771=>x"00037",
772=>x"00037",
773=>x"00037",
774=>x"00037",
775=>x"00037",
776=>x"00037",
777=>x"00037",
778=>x"00037",
779=>x"00037",
780=>x"00037",
781=>x"00037",
782=>x"00037",
783=>x"00037",
784=>x"00038",
785=>x"00038",
786=>x"00038",
787=>x"00038",
788=>x"00038",
789=>x"00038",
790=>x"00038",
791=>x"00038",
792=>x"00038",
793=>x"00038",
794=>x"00038",
795=>x"00038",
796=>x"00038",
797=>x"00038",
798=>x"00039",
799=>x"00039",
800=>x"00039",
801=>x"00039",
802=>x"00039",
803=>x"00039",
804=>x"00039",
805=>x"00039",
806=>x"00039",
807=>x"00039",
808=>x"00039",
809=>x"00039",
810=>x"00039",
811=>x"00039",
812=>x"0003a",
813=>x"0003a",
814=>x"0003a",
815=>x"0003a",
816=>x"0003a",
817=>x"0003a",
818=>x"0003a",
819=>x"0003a",
820=>x"0003a",
821=>x"0003a",
822=>x"0003a",
823=>x"0003a",
824=>x"0003a",
825=>x"0003a",
826=>x"0003b",
827=>x"0003b",
828=>x"0003b",
829=>x"0003b",
830=>x"0003b",
831=>x"0003b",
832=>x"0003b",
833=>x"0003b",
834=>x"0003b",
835=>x"0003b",
836=>x"0003b",
837=>x"0003b",
838=>x"0003b",
839=>x"0003b",
840=>x"0003c",
841=>x"0003c",
842=>x"0003c",
843=>x"0003c",
844=>x"0003c",
845=>x"0003c",
846=>x"0003c",
847=>x"0003c",
848=>x"0003c",
849=>x"0003c",
850=>x"0003c",
851=>x"0003c",
852=>x"0003c",
853=>x"0003c",
854=>x"0003d",
855=>x"0003d",
856=>x"0003d",
857=>x"0003d",
858=>x"0003d",
859=>x"0003d",
860=>x"0003d",
861=>x"0003d",
862=>x"0003d",
863=>x"0003d",
864=>x"0003d",
865=>x"0003d",
866=>x"0003d",
867=>x"0003d",
868=>x"0003e",
869=>x"0003e",
870=>x"0003e",
871=>x"0003e",
872=>x"0003e",
873=>x"0003e",
874=>x"0003e",
875=>x"0003e",
876=>x"0003e",
877=>x"0003e",
878=>x"0003e",
879=>x"0003e",
880=>x"0003e",
881=>x"0003e",
882=>x"0003f",
883=>x"0003f",
884=>x"0003f",
885=>x"0003f",
886=>x"0003f",
887=>x"0003f",
888=>x"0003f",
889=>x"0003f",
890=>x"0003f",
891=>x"0003f",
892=>x"0003f",
893=>x"0003f",
894=>x"0003f",
895=>x"0003f",
896=>x"00040",
897=>x"00040",
898=>x"00040",
899=>x"00040",
900=>x"00040",
901=>x"00040",
902=>x"00040",
903=>x"00040",
904=>x"00040",
905=>x"00040",
906=>x"00040",
907=>x"00040",
908=>x"00040",
909=>x"00040",
910=>x"00041",
911=>x"00041",
912=>x"00041",
913=>x"00041",
914=>x"00041",
915=>x"00041",
916=>x"00041",
917=>x"00041",
918=>x"00041",
919=>x"00041",
920=>x"00041",
921=>x"00041",
922=>x"00041",
923=>x"00041",
924=>x"00042",
925=>x"00042",
926=>x"00042",
927=>x"00042",
928=>x"00042",
929=>x"00042",
930=>x"00042",
931=>x"00042",
932=>x"00042",
933=>x"00042",
934=>x"00042",
935=>x"00042",
936=>x"00042",
937=>x"00042",
938=>x"00043",
939=>x"00043",
940=>x"00043",
941=>x"00043",
942=>x"00043",
943=>x"00043",
944=>x"00043",
945=>x"00043",
946=>x"00043",
947=>x"00043",
948=>x"00043",
949=>x"00043",
950=>x"00043",
951=>x"00043",
952=>x"00044",
953=>x"00044",
954=>x"00044",
955=>x"00044",
956=>x"00044",
957=>x"00044",
958=>x"00044",
959=>x"00044",
960=>x"00044",
961=>x"00044",
962=>x"00044",
963=>x"00044",
964=>x"00044",
965=>x"00044",
966=>x"00045",
967=>x"00045",
968=>x"00045",
969=>x"00045",
970=>x"00045",
971=>x"00045",
972=>x"00045",
973=>x"00045",
974=>x"00045",
975=>x"00045",
976=>x"00045",
977=>x"00045",
978=>x"00045",
979=>x"00045",
980=>x"00046",
981=>x"00046",
982=>x"00046",
983=>x"00046",
984=>x"00046",
985=>x"00046",
986=>x"00046",
987=>x"00046",
988=>x"00046",
989=>x"00046",
990=>x"00046",
991=>x"00046",
992=>x"00046",
993=>x"00046",
994=>x"00047",
995=>x"00047",
996=>x"00047",
997=>x"00047",
998=>x"00047",
999=>x"00047",
1000=>x"00047",
1001=>x"00047",
1002=>x"00047",
1003=>x"00047",
1004=>x"00047",
1005=>x"00047",
1006=>x"00047",
1007=>x"00047",
1008=>x"00048",
1009=>x"00048",
1010=>x"00048",
1011=>x"00048",
1012=>x"00048",
1013=>x"00048",
1014=>x"00048",
1015=>x"00048",
1016=>x"00048",
1017=>x"00048",
1018=>x"00048",
1019=>x"00048",
1020=>x"00048",
1021=>x"00048",
1022=>x"00049",
1023=>x"00049",
1024=>x"00049",
1025=>x"00049",
1026=>x"00049",
1027=>x"00049",
1028=>x"00049",
1029=>x"00049",
1030=>x"00049",
1031=>x"00049",
1032=>x"00049",
1033=>x"00049",
1034=>x"00049",
1035=>x"00049",
1036=>x"0004a",
1037=>x"0004a",
1038=>x"0004a",
1039=>x"0004a",
1040=>x"0004a",
1041=>x"0004a",
1042=>x"0004a",
1043=>x"0004a",
1044=>x"0004a",
1045=>x"0004a",
1046=>x"0004a",
1047=>x"0004a",
1048=>x"0004a",
1049=>x"0004a",
1050=>x"0004b",
1051=>x"0004b",
1052=>x"0004b",
1053=>x"0004b",
1054=>x"0004b",
1055=>x"0004b",
1056=>x"0004b",
1057=>x"0004b",
1058=>x"0004b",
1059=>x"0004b",
1060=>x"0004b",
1061=>x"0004b",
1062=>x"0004b",
1063=>x"0004b",
1064=>x"0004c",
1065=>x"0004c",
1066=>x"0004c",
1067=>x"0004c",
1068=>x"0004c",
1069=>x"0004c",
1070=>x"0004c",
1071=>x"0004c",
1072=>x"0004c",
1073=>x"0004c",
1074=>x"0004c",
1075=>x"0004c",
1076=>x"0004c",
1077=>x"0004c",
1078=>x"0004d",
1079=>x"0004d",
1080=>x"0004d",
1081=>x"0004d",
1082=>x"0004d",
1083=>x"0004d",
1084=>x"0004d",
1085=>x"0004d",
1086=>x"0004d",
1087=>x"0004d",
1088=>x"0004d",
1089=>x"0004d",
1090=>x"0004d",
1091=>x"0004d",
1092=>x"0004e",
1093=>x"0004e",
1094=>x"0004e",
1095=>x"0004e",
1096=>x"0004e",
1097=>x"0004e",
1098=>x"0004e",
1099=>x"0004e",
1100=>x"0004e",
1101=>x"0004e",
1102=>x"0004e",
1103=>x"0004e",
1104=>x"0004e",
1105=>x"0004e",
1106=>x"0004f",
1107=>x"0004f",
1108=>x"0004f",
1109=>x"0004f",
1110=>x"0004f",
1111=>x"0004f",
1112=>x"0004f",
1113=>x"0004f",
1114=>x"0004f",
1115=>x"0004f",
1116=>x"0004f",
1117=>x"0004f",
1118=>x"0004f",
1119=>x"0004f",
1120=>x"00050",
1121=>x"00050",
1122=>x"00050",
1123=>x"00050",
1124=>x"00050",
1125=>x"00050",
1126=>x"00050",
1127=>x"00050",
1128=>x"00050",
1129=>x"00050",
1130=>x"00050",
1131=>x"00050",
1132=>x"00050",
1133=>x"00050",
1134=>x"00051",
1135=>x"00051",
1136=>x"00051",
1137=>x"00051",
1138=>x"00051",
1139=>x"00051",
1140=>x"00051",
1141=>x"00051",
1142=>x"00051",
1143=>x"00051",
1144=>x"00051",
1145=>x"00051",
1146=>x"00051",
1147=>x"00051",
1148=>x"00052",
1149=>x"00052",
1150=>x"00052",
1151=>x"00052",
1152=>x"00052",
1153=>x"00052",
1154=>x"00052",
1155=>x"00052",
1156=>x"00052",
1157=>x"00052",
1158=>x"00052",
1159=>x"00052",
1160=>x"00052",
1161=>x"00052",
1162=>x"00053",
1163=>x"00053",
1164=>x"00053",
1165=>x"00053",
1166=>x"00053",
1167=>x"00053",
1168=>x"00053",
1169=>x"00053",
1170=>x"00053",
1171=>x"00053",
1172=>x"00053",
1173=>x"00053",
1174=>x"00053",
1175=>x"00053",
1176=>x"00054",
1177=>x"00054",
1178=>x"00054",
1179=>x"00054",
1180=>x"00054",
1181=>x"00054",
1182=>x"00054",
1183=>x"00054",
1184=>x"00054",
1185=>x"00054",
1186=>x"00054",
1187=>x"00054",
1188=>x"00054",
1189=>x"00054",
1190=>x"00055",
1191=>x"00055",
1192=>x"00055",
1193=>x"00055",
1194=>x"00055",
1195=>x"00055",
1196=>x"00055",
1197=>x"00055",
1198=>x"00055",
1199=>x"00055",
1200=>x"00055",
1201=>x"00055",
1202=>x"00055",
1203=>x"00055",
1204=>x"00056",
1205=>x"00056",
1206=>x"00056",
1207=>x"00056",
1208=>x"00056",
1209=>x"00056",
1210=>x"00056",
1211=>x"00056",
1212=>x"00056",
1213=>x"00056",
1214=>x"00056",
1215=>x"00056",
1216=>x"00056",
1217=>x"00056",
1218=>x"00057",
1219=>x"00057",
1220=>x"00057",
1221=>x"00057",
1222=>x"00057",
1223=>x"00057",
1224=>x"00057",
1225=>x"00057",
1226=>x"00057",
1227=>x"00057",
1228=>x"00057",
1229=>x"00057",
1230=>x"00057",
1231=>x"00057",
1232=>x"00058",
1233=>x"00058",
1234=>x"00058",
1235=>x"00058",
1236=>x"00058",
1237=>x"00058",
1238=>x"00058",
1239=>x"00058",
1240=>x"00058",
1241=>x"00058",
1242=>x"00058",
1243=>x"00058",
1244=>x"00058",
1245=>x"00058",
1246=>x"00059",
1247=>x"00059",
1248=>x"00059",
1249=>x"00059",
1250=>x"00059",
1251=>x"00059",
1252=>x"00059",
1253=>x"00059",
1254=>x"00059",
1255=>x"00059",
1256=>x"00059",
1257=>x"00059",
1258=>x"00059",
1259=>x"00059",
1260=>x"0005a",
1261=>x"0005a",
1262=>x"0005a",
1263=>x"0005a",
1264=>x"0005a",
1265=>x"0005a",
1266=>x"0005a",
1267=>x"0005a",
1268=>x"0005a",
1269=>x"0005a",
1270=>x"0005a",
1271=>x"0005a",
1272=>x"0005a",
1273=>x"0005a",
1274=>x"0005b",
1275=>x"0005b",
1276=>x"0005b",
1277=>x"0005b",
1278=>x"0005b",
1279=>x"0005b",
1280=>x"0005b",
1281=>x"0005b",
1282=>x"0005b",
1283=>x"0005b",
1284=>x"0005b",
1285=>x"0005b",
1286=>x"0005b",
1287=>x"0005b",
1288=>x"0005c",
1289=>x"0005c",
1290=>x"0005c",
1291=>x"0005c",
1292=>x"0005c",
1293=>x"0005c",
1294=>x"0005c",
1295=>x"0005c",
1296=>x"0005c",
1297=>x"0005c",
1298=>x"0005c",
1299=>x"0005c",
1300=>x"0005c",
1301=>x"0005c",
1302=>x"0005d",
1303=>x"0005d",
1304=>x"0005d",
1305=>x"0005d",
1306=>x"0005d",
1307=>x"0005d",
1308=>x"0005d",
1309=>x"0005d",
1310=>x"0005d",
1311=>x"0005d",
1312=>x"0005d",
1313=>x"0005d",
1314=>x"0005d",
1315=>x"0005d",
1316=>x"0005e",
1317=>x"0005e",
1318=>x"0005e",
1319=>x"0005e",
1320=>x"0005e",
1321=>x"0005e",
1322=>x"0005e",
1323=>x"0005e",
1324=>x"0005e",
1325=>x"0005e",
1326=>x"0005e",
1327=>x"0005e",
1328=>x"0005e",
1329=>x"0005e",
1330=>x"0005f",
1331=>x"0005f",
1332=>x"0005f",
1333=>x"0005f",
1334=>x"0005f",
1335=>x"0005f",
1336=>x"0005f",
1337=>x"0005f",
1338=>x"0005f",
1339=>x"0005f",
1340=>x"0005f",
1341=>x"0005f",
1342=>x"0005f",
1343=>x"0005f",
1344=>x"00060",
1345=>x"00060",
1346=>x"00060",
1347=>x"00060",
1348=>x"00060",
1349=>x"00060",
1350=>x"00060",
1351=>x"00060",
1352=>x"00060",
1353=>x"00060",
1354=>x"00060",
1355=>x"00060",
1356=>x"00060",
1357=>x"00060",
1358=>x"00061",
1359=>x"00061",
1360=>x"00061",
1361=>x"00061",
1362=>x"00061",
1363=>x"00061",
1364=>x"00061",
1365=>x"00061",
1366=>x"00061",
1367=>x"00061",
1368=>x"00061",
1369=>x"00061",
1370=>x"00061",
1371=>x"00061",
1372=>x"00062",
1373=>x"00062",
1374=>x"00062",
1375=>x"00062",
1376=>x"00062",
1377=>x"00062",
1378=>x"00062",
1379=>x"00062",
1380=>x"00062",
1381=>x"00062",
1382=>x"00062",
1383=>x"00062",
1384=>x"00062",
1385=>x"00062",
1386=>x"00063",
1387=>x"00063",
1388=>x"00063",
1389=>x"00063",
1390=>x"00063",
1391=>x"00063",
1392=>x"00063",
1393=>x"00063",
1394=>x"00063",
1395=>x"00063",
1396=>x"00063",
1397=>x"00063",
1398=>x"00063",
1399=>x"00063",
1400=>x"00064",
1401=>x"00064",
1402=>x"00064",
1403=>x"00064",
1404=>x"00064",
1405=>x"00064",
1406=>x"00064",
1407=>x"00064",
1408=>x"00064",
1409=>x"00064",
1410=>x"00064",
1411=>x"00064",
1412=>x"00064",
1413=>x"00064",
1414=>x"00065",
1415=>x"00065",
1416=>x"00065",
1417=>x"00065",
1418=>x"00065",
1419=>x"00065",
1420=>x"00065",
1421=>x"00065",
1422=>x"00065",
1423=>x"00065",
1424=>x"00065",
1425=>x"00065",
1426=>x"00065",
1427=>x"00065",
1428=>x"00066",
1429=>x"00066",
1430=>x"00066",
1431=>x"00066",
1432=>x"00066",
1433=>x"00066",
1434=>x"00066",
1435=>x"00066",
1436=>x"00066",
1437=>x"00066",
1438=>x"00066",
1439=>x"00066",
1440=>x"00066",
1441=>x"00066",
1442=>x"00067",
1443=>x"00067",
1444=>x"00067",
1445=>x"00067",
1446=>x"00067",
1447=>x"00067",
1448=>x"00067",
1449=>x"00067",
1450=>x"00067",
1451=>x"00067",
1452=>x"00067",
1453=>x"00067",
1454=>x"00067",
1455=>x"00067",
1456=>x"00068",
1457=>x"00068",
1458=>x"00068",
1459=>x"00068",
1460=>x"00068",
1461=>x"00068",
1462=>x"00068",
1463=>x"00068",
1464=>x"00068",
1465=>x"00068",
1466=>x"00068",
1467=>x"00068",
1468=>x"00068",
1469=>x"00068",
1470=>x"00069",
1471=>x"00069",
1472=>x"00069",
1473=>x"00069",
1474=>x"00069",
1475=>x"00069",
1476=>x"00069",
1477=>x"00069",
1478=>x"00069",
1479=>x"00069",
1480=>x"00069",
1481=>x"00069",
1482=>x"00069",
1483=>x"00069",
1484=>x"0006a",
1485=>x"0006a",
1486=>x"0006a",
1487=>x"0006a",
1488=>x"0006a",
1489=>x"0006a",
1490=>x"0006a",
1491=>x"0006a",
1492=>x"0006a",
1493=>x"0006a",
1494=>x"0006a",
1495=>x"0006a",
1496=>x"0006a",
1497=>x"0006a",
1498=>x"0006b",
1499=>x"0006b",
1500=>x"0006b",
1501=>x"0006b",
1502=>x"0006b",
1503=>x"0006b",
1504=>x"0006b",
1505=>x"0006b",
1506=>x"0006b",
1507=>x"0006b",
1508=>x"0006b",
1509=>x"0006b",
1510=>x"0006b",
1511=>x"0006b",
1512=>x"0006c",
1513=>x"0006c",
1514=>x"0006c",
1515=>x"0006c",
1516=>x"0006c",
1517=>x"0006c",
1518=>x"0006c",
1519=>x"0006c",
1520=>x"0006c",
1521=>x"0006c",
1522=>x"0006c",
1523=>x"0006c",
1524=>x"0006c",
1525=>x"0006c",
1526=>x"0006d",
1527=>x"0006d",
1528=>x"0006d",
1529=>x"0006d",
1530=>x"0006d",
1531=>x"0006d",
1532=>x"0006d",
1533=>x"0006d",
1534=>x"0006d",
1535=>x"0006d",
1536=>x"0006d",
1537=>x"0006d",
1538=>x"0006d",
1539=>x"0006d",
1540=>x"0006e",
1541=>x"0006e",
1542=>x"0006e",
1543=>x"0006e",
1544=>x"0006e",
1545=>x"0006e",
1546=>x"0006e",
1547=>x"0006e",
1548=>x"0006e",
1549=>x"0006e",
1550=>x"0006e",
1551=>x"0006e",
1552=>x"0006e",
1553=>x"0006e",
1554=>x"0006f",
1555=>x"0006f",
1556=>x"0006f",
1557=>x"0006f",
1558=>x"0006f",
1559=>x"0006f",
1560=>x"0006f",
1561=>x"0006f",
1562=>x"0006f",
1563=>x"0006f",
1564=>x"0006f",
1565=>x"0006f",
1566=>x"0006f",
1567=>x"0006f",
1568=>x"00070",
1569=>x"00070",
1570=>x"00070",
1571=>x"00070",
1572=>x"00070",
1573=>x"00070",
1574=>x"00070",
1575=>x"00070",
1576=>x"00070",
1577=>x"00070",
1578=>x"00070",
1579=>x"00070",
1580=>x"00070",
1581=>x"00070",
1582=>x"00071",
1583=>x"00071",
1584=>x"00071",
1585=>x"00071",
1586=>x"00071",
1587=>x"00071",
1588=>x"00071",
1589=>x"00071",
1590=>x"00071",
1591=>x"00071",
1592=>x"00071",
1593=>x"00071",
1594=>x"00071",
1595=>x"00071",
1596=>x"00072",
1597=>x"00072",
1598=>x"00072",
1599=>x"00072",
1600=>x"00072",
1601=>x"00072",
1602=>x"00072",
1603=>x"00072",
1604=>x"00072",
1605=>x"00072",
1606=>x"00072",
1607=>x"00072",
1608=>x"00072",
1609=>x"00072",
1610=>x"00073",
1611=>x"00073",
1612=>x"00073",
1613=>x"00073",
1614=>x"00073",
1615=>x"00073",
1616=>x"00073",
1617=>x"00073",
1618=>x"00073",
1619=>x"00073",
1620=>x"00073",
1621=>x"00073",
1622=>x"00073",
1623=>x"00073",
1624=>x"00074",
1625=>x"00074",
1626=>x"00074",
1627=>x"00074",
1628=>x"00074",
1629=>x"00074",
1630=>x"00074",
1631=>x"00074",
1632=>x"00074",
1633=>x"00074",
1634=>x"00074",
1635=>x"00074",
1636=>x"00074",
1637=>x"00074",
1638=>x"00075",
1639=>x"00075",
1640=>x"00075",
1641=>x"00075",
1642=>x"00075",
1643=>x"00075",
1644=>x"00075",
1645=>x"00075",
1646=>x"00075",
1647=>x"00075",
1648=>x"00075",
1649=>x"00075",
1650=>x"00075",
1651=>x"00075",
1652=>x"00076",
1653=>x"00076",
1654=>x"00076",
1655=>x"00076",
1656=>x"00076",
1657=>x"00076",
1658=>x"00076",
1659=>x"00076",
1660=>x"00076",
1661=>x"00076",
1662=>x"00076",
1663=>x"00076",
1664=>x"00076",
1665=>x"00076",
1666=>x"00077",
1667=>x"00077",
1668=>x"00077",
1669=>x"00077",
1670=>x"00077",
1671=>x"00077",
1672=>x"00077",
1673=>x"00077",
1674=>x"00077",
1675=>x"00077",
1676=>x"00077",
1677=>x"00077",
1678=>x"00077",
1679=>x"00077",
1680=>x"00078",
1681=>x"00078",
1682=>x"00078",
1683=>x"00078",
1684=>x"00078",
1685=>x"00078",
1686=>x"00078",
1687=>x"00078",
1688=>x"00078",
1689=>x"00078",
1690=>x"00078",
1691=>x"00078",
1692=>x"00078",
1693=>x"00078",
1694=>x"00079",
1695=>x"00079",
1696=>x"00079",
1697=>x"00079",
1698=>x"00079",
1699=>x"00079",
1700=>x"00079",
1701=>x"00079",
1702=>x"00079",
1703=>x"00079",
1704=>x"00079",
1705=>x"00079",
1706=>x"00079",
1707=>x"00079",
1708=>x"0007a",
1709=>x"0007a",
1710=>x"0007a",
1711=>x"0007a",
1712=>x"0007a",
1713=>x"0007a",
1714=>x"0007a",
1715=>x"0007a",
1716=>x"0007a",
1717=>x"0007a",
1718=>x"0007a",
1719=>x"0007a",
1720=>x"0007a",
1721=>x"0007a",
1722=>x"0007b",
1723=>x"0007b",
1724=>x"0007b",
1725=>x"0007b",
1726=>x"0007b",
1727=>x"0007b",
1728=>x"0007b",
1729=>x"0007b",
1730=>x"0007b",
1731=>x"0007b",
1732=>x"0007b",
1733=>x"0007b",
1734=>x"0007b",
1735=>x"0007b",
1736=>x"0007c",
1737=>x"0007c",
1738=>x"0007c",
1739=>x"0007c",
1740=>x"0007c",
1741=>x"0007c",
1742=>x"0007c",
1743=>x"0007c",
1744=>x"0007c",
1745=>x"0007c",
1746=>x"0007c",
1747=>x"0007c",
1748=>x"0007c",
1749=>x"0007c",
1750=>x"0007d",
1751=>x"0007d",
1752=>x"0007d",
1753=>x"0007d",
1754=>x"0007d",
1755=>x"0007d",
1756=>x"0007d",
1757=>x"0007d",
1758=>x"0007d",
1759=>x"0007d",
1760=>x"0007d",
1761=>x"0007d",
1762=>x"0007d",
1763=>x"0007d",
1764=>x"0007e",
1765=>x"0007e",
1766=>x"0007e",
1767=>x"0007e",
1768=>x"0007e",
1769=>x"0007e",
1770=>x"0007e",
1771=>x"0007e",
1772=>x"0007e",
1773=>x"0007e",
1774=>x"0007e",
1775=>x"0007e",
1776=>x"0007e",
1777=>x"0007e",
1778=>x"0007f",
1779=>x"0007f",
1780=>x"0007f",
1781=>x"0007f",
1782=>x"0007f",
1783=>x"0007f",
1784=>x"0007f",
1785=>x"0007f",
1786=>x"0007f",
1787=>x"0007f",
1788=>x"0007f",
1789=>x"0007f",
1790=>x"0007f",
1791=>x"0007f",
1792=>x"00080",
1793=>x"00080",
1794=>x"00080",
1795=>x"00080",
1796=>x"00080",
1797=>x"00080",
1798=>x"00080",
1799=>x"00080",
1800=>x"00080",
1801=>x"00080",
1802=>x"00080",
1803=>x"00080",
1804=>x"00080",
1805=>x"00080",
1806=>x"00081",
1807=>x"00081",
1808=>x"00081",
1809=>x"00081",
1810=>x"00081",
1811=>x"00081",
1812=>x"00081",
1813=>x"00081",
1814=>x"00081",
1815=>x"00081",
1816=>x"00081",
1817=>x"00081",
1818=>x"00081",
1819=>x"00081",
1820=>x"00082",
1821=>x"00082",
1822=>x"00082",
1823=>x"00082",
1824=>x"00082",
1825=>x"00082",
1826=>x"00082",
1827=>x"00082",
1828=>x"00082",
1829=>x"00082",
1830=>x"00082",
1831=>x"00082",
1832=>x"00082",
1833=>x"00082",
1834=>x"00083",
1835=>x"00083",
1836=>x"00083",
1837=>x"00083",
1838=>x"00083",
1839=>x"00083",
1840=>x"00083",
1841=>x"00083",
1842=>x"00083",
1843=>x"00083",
1844=>x"00083",
1845=>x"00083",
1846=>x"00083",
1847=>x"00083",
1848=>x"00084",
1849=>x"00084",
1850=>x"00084",
1851=>x"00084",
1852=>x"00084",
1853=>x"00084",
1854=>x"00084",
1855=>x"00084",
1856=>x"00084",
1857=>x"00084",
1858=>x"00084",
1859=>x"00084",
1860=>x"00084",
1861=>x"00084",
1862=>x"00085",
1863=>x"00085",
1864=>x"00085",
1865=>x"00085",
1866=>x"00085",
1867=>x"00085",
1868=>x"00085",
1869=>x"00085",
1870=>x"00085",
1871=>x"00085",
1872=>x"00085",
1873=>x"00085",
1874=>x"00085",
1875=>x"00085",
1876=>x"00086",
1877=>x"00086",
1878=>x"00086",
1879=>x"00086",
1880=>x"00086",
1881=>x"00086",
1882=>x"00086",
1883=>x"00086",
1884=>x"00086",
1885=>x"00086",
1886=>x"00086",
1887=>x"00086",
1888=>x"00086",
1889=>x"00086",
1890=>x"00087",
1891=>x"00087",
1892=>x"00087",
1893=>x"00087",
1894=>x"00087",
1895=>x"00087",
1896=>x"00087",
1897=>x"00087",
1898=>x"00087",
1899=>x"00087",
1900=>x"00087",
1901=>x"00087",
1902=>x"00087",
1903=>x"00087",
1904=>x"00088",
1905=>x"00088",
1906=>x"00088",
1907=>x"00088",
1908=>x"00088",
1909=>x"00088",
1910=>x"00088",
1911=>x"00088",
1912=>x"00088",
1913=>x"00088",
1914=>x"00088",
1915=>x"00088",
1916=>x"00088",
1917=>x"00088",
1918=>x"00089",
1919=>x"00089",
1920=>x"00089",
1921=>x"00089",
1922=>x"00089",
1923=>x"00089",
1924=>x"00089",
1925=>x"00089",
1926=>x"00089",
1927=>x"00089",
1928=>x"00089",
1929=>x"00089",
1930=>x"00089",
1931=>x"00089",
1932=>x"0008a",
1933=>x"0008a",
1934=>x"0008a",
1935=>x"0008a",
1936=>x"0008a",
1937=>x"0008a",
1938=>x"0008a",
1939=>x"0008a",
1940=>x"0008a",
1941=>x"0008a",
1942=>x"0008a",
1943=>x"0008a",
1944=>x"0008a",
1945=>x"0008a",
1946=>x"0008b",
1947=>x"0008b",
1948=>x"0008b",
1949=>x"0008b",
1950=>x"0008b",
1951=>x"0008b",
1952=>x"0008b",
1953=>x"0008b",
1954=>x"0008b",
1955=>x"0008b",
1956=>x"0008b",
1957=>x"0008b",
1958=>x"0008b",
1959=>x"0008b",
1960=>x"0008c",
1961=>x"0008c",
1962=>x"0008c",
1963=>x"0008c",
1964=>x"0008c",
1965=>x"0008c",
1966=>x"0008c",
1967=>x"0008c",
1968=>x"0008c",
1969=>x"0008c",
1970=>x"0008c",
1971=>x"0008c",
1972=>x"0008c",
1973=>x"0008c",
1974=>x"0008d",
1975=>x"0008d",
1976=>x"0008d",
1977=>x"0008d",
1978=>x"0008d",
1979=>x"0008d",
1980=>x"0008d",
1981=>x"0008d",
1982=>x"0008d",
1983=>x"0008d",
1984=>x"0008d",
1985=>x"0008d",
1986=>x"0008d",
1987=>x"0008d",
1988=>x"0008e",
1989=>x"0008e",
1990=>x"0008e",
1991=>x"0008e",
1992=>x"0008e",
1993=>x"0008e",
1994=>x"0008e",
1995=>x"0008e",
1996=>x"0008e",
1997=>x"0008e",
1998=>x"0008e",
1999=>x"0008e",
2000=>x"0008e",
2001=>x"0008e",
2002=>x"0008f",
2003=>x"0008f",
2004=>x"0008f",
2005=>x"0008f",
2006=>x"0008f",
2007=>x"0008f",
2008=>x"0008f",
2009=>x"0008f",
2010=>x"0008f",
2011=>x"0008f",
2012=>x"0008f",
2013=>x"0008f",
2014=>x"0008f",
2015=>x"0008f",
2016=>x"00090",
2017=>x"00090",
2018=>x"00090",
2019=>x"00090",
2020=>x"00090",
2021=>x"00090",
2022=>x"00090",
2023=>x"00090",
2024=>x"00090",
2025=>x"00090",
2026=>x"00090",
2027=>x"00090",
2028=>x"00090",
2029=>x"00090",
2030=>x"00091",
2031=>x"00091",
2032=>x"00091",
2033=>x"00091",
2034=>x"00091",
2035=>x"00091",
2036=>x"00091",
2037=>x"00091",
2038=>x"00091",
2039=>x"00091",
2040=>x"00091",
2041=>x"00091",
2042=>x"00091",
2043=>x"00091",
2044=>x"00092",
2045=>x"00092",
2046=>x"00092",
2047=>x"00092",
2048=>x"00092",
2049=>x"00092",
2050=>x"00092",
2051=>x"00092",
2052=>x"00092",
2053=>x"00092",
2054=>x"00092",
2055=>x"00092",
2056=>x"00092",
2057=>x"00092",
2058=>x"00093",
2059=>x"00093",
2060=>x"00093",
2061=>x"00093",
2062=>x"00093",
2063=>x"00093",
2064=>x"00093",
2065=>x"00093",
2066=>x"00093",
2067=>x"00093",
2068=>x"00093",
2069=>x"00093",
2070=>x"00093",
2071=>x"00093",
2072=>x"00094",
2073=>x"00094",
2074=>x"00094",
2075=>x"00094",
2076=>x"00094",
2077=>x"00094",
2078=>x"00094",
2079=>x"00094",
2080=>x"00094",
2081=>x"00094",
2082=>x"00094",
2083=>x"00094",
2084=>x"00094",
2085=>x"00094",
2086=>x"00095",
2087=>x"00095",
2088=>x"00095",
2089=>x"00095",
2090=>x"00095",
2091=>x"00095",
2092=>x"00095",
2093=>x"00095",
2094=>x"00095",
2095=>x"00095",
2096=>x"00095",
2097=>x"00095",
2098=>x"00095",
2099=>x"00095",
2100=>x"00096",
2101=>x"00096",
2102=>x"00096",
2103=>x"00096",
2104=>x"00096",
2105=>x"00096",
2106=>x"00096",
2107=>x"00096",
2108=>x"00096",
2109=>x"00096",
2110=>x"00096",
2111=>x"00096",
2112=>x"00096",
2113=>x"00096",
2114=>x"00097",
2115=>x"00097",
2116=>x"00097",
2117=>x"00097",
2118=>x"00097",
2119=>x"00097",
2120=>x"00097",
2121=>x"00097",
2122=>x"00097",
2123=>x"00097",
2124=>x"00097",
2125=>x"00097",
2126=>x"00097",
2127=>x"00097",
2128=>x"00098",
2129=>x"00098",
2130=>x"00098",
2131=>x"00098",
2132=>x"00098",
2133=>x"00098",
2134=>x"00098",
2135=>x"00098",
2136=>x"00098",
2137=>x"00098",
2138=>x"00098",
2139=>x"00098",
2140=>x"00098",
2141=>x"00098",
2142=>x"00099",
2143=>x"00099",
2144=>x"00099",
2145=>x"00099",
2146=>x"00099",
2147=>x"00099",
2148=>x"00099",
2149=>x"00099",
2150=>x"00099",
2151=>x"00099",
2152=>x"00099",
2153=>x"00099",
2154=>x"00099",
2155=>x"00099",
2156=>x"0009a",
2157=>x"0009a",
2158=>x"0009a",
2159=>x"0009a",
2160=>x"0009a",
2161=>x"0009a",
2162=>x"0009a",
2163=>x"0009a",
2164=>x"0009a",
2165=>x"0009a",
2166=>x"0009a",
2167=>x"0009a",
2168=>x"0009a",
2169=>x"0009a",
2170=>x"0009b",
2171=>x"0009b",
2172=>x"0009b",
2173=>x"0009b",
2174=>x"0009b",
2175=>x"0009b",
2176=>x"0009b",
2177=>x"0009b",
2178=>x"0009b",
2179=>x"0009b",
2180=>x"0009b",
2181=>x"0009b",
2182=>x"0009b",
2183=>x"0009b",
2184=>x"0009c",
2185=>x"0009c",
2186=>x"0009c",
2187=>x"0009c",
2188=>x"0009c",
2189=>x"0009c",
2190=>x"0009c",
2191=>x"0009c",
2192=>x"0009c",
2193=>x"0009c",
2194=>x"0009c",
2195=>x"0009c",
2196=>x"0009c",
2197=>x"0009c",
2198=>x"0009d",
2199=>x"0009d",
2200=>x"0009d",
2201=>x"0009d",
2202=>x"0009d",
2203=>x"0009d",
2204=>x"0009d",
2205=>x"0009d",
2206=>x"0009d",
2207=>x"0009d",
2208=>x"0009d",
2209=>x"0009d",
2210=>x"0009d",
2211=>x"0009d",
2212=>x"0009e",
2213=>x"0009e",
2214=>x"0009e",
2215=>x"0009e",
2216=>x"0009e",
2217=>x"0009e",
2218=>x"0009e",
2219=>x"0009e",
2220=>x"0009e",
2221=>x"0009e",
2222=>x"0009e",
2223=>x"0009e",
2224=>x"0009e",
2225=>x"0009e",
2226=>x"0009f",
2227=>x"0009f",
2228=>x"0009f",
2229=>x"0009f",
2230=>x"0009f",
2231=>x"0009f",
2232=>x"0009f",
2233=>x"0009f",
2234=>x"0009f",
2235=>x"0009f",
2236=>x"0009f",
2237=>x"0009f",
2238=>x"0009f",
2239=>x"0009f",
2240=>x"000a0",
2241=>x"000a0",
2242=>x"000a0",
2243=>x"000a0",
2244=>x"000a0",
2245=>x"000a0",
2246=>x"000a0",
2247=>x"000a0",
2248=>x"000a0",
2249=>x"000a0",
2250=>x"000a0",
2251=>x"000a0",
2252=>x"000a0",
2253=>x"000a0",
2254=>x"000a1",
2255=>x"000a1",
2256=>x"000a1",
2257=>x"000a1",
2258=>x"000a1",
2259=>x"000a1",
2260=>x"000a1",
2261=>x"000a1",
2262=>x"000a1",
2263=>x"000a1",
2264=>x"000a1",
2265=>x"000a1",
2266=>x"000a1",
2267=>x"000a1",
2268=>x"000a2",
2269=>x"000a2",
2270=>x"000a2",
2271=>x"000a2",
2272=>x"000a2",
2273=>x"000a2",
2274=>x"000a2",
2275=>x"000a2",
2276=>x"000a2",
2277=>x"000a2",
2278=>x"000a2",
2279=>x"000a2",
2280=>x"000a2",
2281=>x"000a2",
2282=>x"000a3",
2283=>x"000a3",
2284=>x"000a3",
2285=>x"000a3",
2286=>x"000a3",
2287=>x"000a3",
2288=>x"000a3",
2289=>x"000a3",
2290=>x"000a3",
2291=>x"000a3",
2292=>x"000a3",
2293=>x"000a3",
2294=>x"000a3",
2295=>x"000a3",
2296=>x"000a4",
2297=>x"000a4",
2298=>x"000a4",
2299=>x"000a4",
2300=>x"000a4",
2301=>x"000a4",
2302=>x"000a4",
2303=>x"000a4",
2304=>x"000a4",
2305=>x"000a4",
2306=>x"000a4",
2307=>x"000a4",
2308=>x"000a4",
2309=>x"000a4",
2310=>x"000a5",
2311=>x"000a5",
2312=>x"000a5",
2313=>x"000a5",
2314=>x"000a5",
2315=>x"000a5",
2316=>x"000a5",
2317=>x"000a5",
2318=>x"000a5",
2319=>x"000a5",
2320=>x"000a5",
2321=>x"000a5",
2322=>x"000a5",
2323=>x"000a5",
2324=>x"000a6",
2325=>x"000a6",
2326=>x"000a6",
2327=>x"000a6",
2328=>x"000a6",
2329=>x"000a6",
2330=>x"000a6",
2331=>x"000a6",
2332=>x"000a6",
2333=>x"000a6",
2334=>x"000a6",
2335=>x"000a6",
2336=>x"000a6",
2337=>x"000a6",
2338=>x"000a7",
2339=>x"000a7",
2340=>x"000a7",
2341=>x"000a7",
2342=>x"000a7",
2343=>x"000a7",
2344=>x"000a7",
2345=>x"000a7",
2346=>x"000a7",
2347=>x"000a7",
2348=>x"000a7",
2349=>x"000a7",
2350=>x"000a7",
2351=>x"000a7",
2352=>x"000a8",
2353=>x"000a8",
2354=>x"000a8",
2355=>x"000a8",
2356=>x"000a8",
2357=>x"000a8",
2358=>x"000a8",
2359=>x"000a8",
2360=>x"000a8",
2361=>x"000a8",
2362=>x"000a8",
2363=>x"000a8",
2364=>x"000a8",
2365=>x"000a8",
2366=>x"000a9",
2367=>x"000a9",
2368=>x"000a9",
2369=>x"000a9",
2370=>x"000a9",
2371=>x"000a9",
2372=>x"000a9",
2373=>x"000a9",
2374=>x"000a9",
2375=>x"000a9",
2376=>x"000a9",
2377=>x"000a9",
2378=>x"000a9",
2379=>x"000a9",
2380=>x"000aa",
2381=>x"000aa",
2382=>x"000aa",
2383=>x"000aa",
2384=>x"000aa",
2385=>x"000aa",
2386=>x"000aa",
2387=>x"000aa",
2388=>x"000aa",
2389=>x"000aa",
2390=>x"000aa",
2391=>x"000aa",
2392=>x"000aa",
2393=>x"000aa",
2394=>x"000ab",
2395=>x"000ab",
2396=>x"000ab",
2397=>x"000ab",
2398=>x"000ab",
2399=>x"000ab",
2400=>x"000ab",
2401=>x"000ab",
2402=>x"000ab",
2403=>x"000ab",
2404=>x"000ab",
2405=>x"000ab",
2406=>x"000ab",
2407=>x"000ab",
2408=>x"000ac",
2409=>x"000ac",
2410=>x"000ac",
2411=>x"000ac",
2412=>x"000ac",
2413=>x"000ac",
2414=>x"000ac",
2415=>x"000ac",
2416=>x"000ac",
2417=>x"000ac",
2418=>x"000ac",
2419=>x"000ac",
2420=>x"000ac",
2421=>x"000ac",
2422=>x"000ad",
2423=>x"000ad",
2424=>x"000ad",
2425=>x"000ad",
2426=>x"000ad",
2427=>x"000ad",
2428=>x"000ad",
2429=>x"000ad",
2430=>x"000ad",
2431=>x"000ad",
2432=>x"000ad",
2433=>x"000ad",
2434=>x"000ad",
2435=>x"000ad",
2436=>x"000ae",
2437=>x"000ae",
2438=>x"000ae",
2439=>x"000ae",
2440=>x"000ae",
2441=>x"000ae",
2442=>x"000ae",
2443=>x"000ae",
2444=>x"000ae",
2445=>x"000ae",
2446=>x"000ae",
2447=>x"000ae",
2448=>x"000ae",
2449=>x"000ae",
2450=>x"000af",
2451=>x"000af",
2452=>x"000af",
2453=>x"000af",
2454=>x"000af",
2455=>x"000af",
2456=>x"000af",
2457=>x"000af",
2458=>x"000af",
2459=>x"000af",
2460=>x"000af",
2461=>x"000af",
2462=>x"000af",
2463=>x"000af",
2464=>x"000b0",
2465=>x"000b0",
2466=>x"000b0",
2467=>x"000b0",
2468=>x"000b0",
2469=>x"000b0",
2470=>x"000b0",
2471=>x"000b0",
2472=>x"000b0",
2473=>x"000b0",
2474=>x"000b0",
2475=>x"000b0",
2476=>x"000b0",
2477=>x"000b0",
2478=>x"000b1",
2479=>x"000b1",
2480=>x"000b1",
2481=>x"000b1",
2482=>x"000b1",
2483=>x"000b1",
2484=>x"000b1",
2485=>x"000b1",
2486=>x"000b1",
2487=>x"000b1",
2488=>x"000b1",
2489=>x"000b1",
2490=>x"000b1",
2491=>x"000b1",
2492=>x"000b2",
2493=>x"000b2",
2494=>x"000b2",
2495=>x"000b2",
2496=>x"000b2",
2497=>x"000b2",
2498=>x"000b2",
2499=>x"000b2",
2500=>x"000b2",
2501=>x"000b2",
2502=>x"000b2",
2503=>x"000b2",
2504=>x"000b2",
2505=>x"000b2",
2506=>x"000b3",
2507=>x"000b3",
2508=>x"000b3",
2509=>x"000b3",
2510=>x"000b3",
2511=>x"000b3",
2512=>x"000b3",
2513=>x"000b3",
2514=>x"000b3",
2515=>x"000b3",
2516=>x"000b3",
2517=>x"000b3",
2518=>x"000b3",
2519=>x"000b3",
2520=>x"000b4",
2521=>x"000b4",
2522=>x"000b4",
2523=>x"000b4",
2524=>x"000b4",
2525=>x"000b4",
2526=>x"000b4",
2527=>x"000b4",
2528=>x"000b4",
2529=>x"000b4",
2530=>x"000b4",
2531=>x"000b4",
2532=>x"000b4",
2533=>x"000b4",
2534=>x"000b5",
2535=>x"000b5",
2536=>x"000b5",
2537=>x"000b5",
2538=>x"000b5",
2539=>x"000b5",
2540=>x"000b5",
2541=>x"000b5",
2542=>x"000b5",
2543=>x"000b5",
2544=>x"000b5",
2545=>x"000b5",
2546=>x"000b5",
2547=>x"000b5",
2548=>x"000b6",
2549=>x"000b6",
2550=>x"000b6",
2551=>x"000b6",
2552=>x"000b6",
2553=>x"000b6",
2554=>x"000b6",
2555=>x"000b6",
2556=>x"000b6",
2557=>x"000b6",
2558=>x"000b6",
2559=>x"000b6",
2560=>x"000b6",
2561=>x"000b6",
2562=>x"000b7",
2563=>x"000b7",
2564=>x"000b7",
2565=>x"000b7",
2566=>x"000b7",
2567=>x"000b7",
2568=>x"000b7",
2569=>x"000b7",
2570=>x"000b7",
2571=>x"000b7",
2572=>x"000b7",
2573=>x"000b7",
2574=>x"000b7",
2575=>x"000b7",
2576=>x"000b8",
2577=>x"000b8",
2578=>x"000b8",
2579=>x"000b8",
2580=>x"000b8",
2581=>x"000b8",
2582=>x"000b8",
2583=>x"000b8",
2584=>x"000b8",
2585=>x"000b8",
2586=>x"000b8",
2587=>x"000b8",
2588=>x"000b8",
2589=>x"000b8",
2590=>x"000b9",
2591=>x"000b9",
2592=>x"000b9",
2593=>x"000b9",
2594=>x"000b9",
2595=>x"000b9",
2596=>x"000b9",
2597=>x"000b9",
2598=>x"000b9",
2599=>x"000b9",
2600=>x"000b9",
2601=>x"000b9",
2602=>x"000b9",
2603=>x"000b9",
2604=>x"000ba",
2605=>x"000ba",
2606=>x"000ba",
2607=>x"000ba",
2608=>x"000ba",
2609=>x"000ba",
2610=>x"000ba",
2611=>x"000ba",
2612=>x"000ba",
2613=>x"000ba",
2614=>x"000ba",
2615=>x"000ba",
2616=>x"000ba",
2617=>x"000ba",
2618=>x"000bb",
2619=>x"000bb",
2620=>x"000bb",
2621=>x"000bb",
2622=>x"000bb",
2623=>x"000bb",
2624=>x"000bb",
2625=>x"000bb",
2626=>x"000bb",
2627=>x"000bb",
2628=>x"000bb",
2629=>x"000bb",
2630=>x"000bb",
2631=>x"000bb",
2632=>x"000bc",
2633=>x"000bc",
2634=>x"000bc",
2635=>x"000bc",
2636=>x"000bc",
2637=>x"000bc",
2638=>x"000bc",
2639=>x"000bc",
2640=>x"000bc",
2641=>x"000bc",
2642=>x"000bc",
2643=>x"000bc",
2644=>x"000bc",
2645=>x"000bc",
2646=>x"000bd",
2647=>x"000bd",
2648=>x"000bd",
2649=>x"000bd",
2650=>x"000bd",
2651=>x"000bd",
2652=>x"000bd",
2653=>x"000bd",
2654=>x"000bd",
2655=>x"000bd",
2656=>x"000bd",
2657=>x"000bd",
2658=>x"000bd",
2659=>x"000bd",
2660=>x"000be",
2661=>x"000be",
2662=>x"000be",
2663=>x"000be",
2664=>x"000be",
2665=>x"000be",
2666=>x"000be",
2667=>x"000be",
2668=>x"000be",
2669=>x"000be",
2670=>x"000be",
2671=>x"000be",
2672=>x"000be",
2673=>x"000be",
2674=>x"000bf",
2675=>x"000bf",
2676=>x"000bf",
2677=>x"000bf",
2678=>x"000bf",
2679=>x"000bf",
2680=>x"000bf",
2681=>x"000bf",
2682=>x"000bf",
2683=>x"000bf",
2684=>x"000bf",
2685=>x"000bf",
2686=>x"000bf",
2687=>x"000bf",
2688=>x"000c0",
2689=>x"000c0",
2690=>x"000c0",
2691=>x"000c0",
2692=>x"000c0",
2693=>x"000c0",
2694=>x"000c0",
2695=>x"000c0",
2696=>x"000c0",
2697=>x"000c0",
2698=>x"000c0",
2699=>x"000c0",
2700=>x"000c0",
2701=>x"000c0",
2702=>x"000c1",
2703=>x"000c1",
2704=>x"000c1",
2705=>x"000c1",
2706=>x"000c1",
2707=>x"000c1",
2708=>x"000c1",
2709=>x"000c1",
2710=>x"000c1",
2711=>x"000c1",
2712=>x"000c1",
2713=>x"000c1",
2714=>x"000c1",
2715=>x"000c1",
2716=>x"000c2",
2717=>x"000c2",
2718=>x"000c2",
2719=>x"000c2",
2720=>x"000c2",
2721=>x"000c2",
2722=>x"000c2",
2723=>x"000c2",
2724=>x"000c2",
2725=>x"000c2",
2726=>x"000c2",
2727=>x"000c2",
2728=>x"000c2",
2729=>x"000c2",
2730=>x"000c3",
2731=>x"000c3",
2732=>x"000c3",
2733=>x"000c3",
2734=>x"000c3",
2735=>x"000c3",
2736=>x"000c3",
2737=>x"000c3",
2738=>x"000c3",
2739=>x"000c3",
2740=>x"000c3",
2741=>x"000c3",
2742=>x"000c3",
2743=>x"000c3",
2744=>x"000c4",
2745=>x"000c4",
2746=>x"000c4",
2747=>x"000c4",
2748=>x"000c4",
2749=>x"000c4",
2750=>x"000c4",
2751=>x"000c4",
2752=>x"000c4",
2753=>x"000c4",
2754=>x"000c4",
2755=>x"000c4",
2756=>x"000c4",
2757=>x"000c4",
2758=>x"000c5",
2759=>x"000c5",
2760=>x"000c5",
2761=>x"000c5",
2762=>x"000c5",
2763=>x"000c5",
2764=>x"000c5",
2765=>x"000c5",
2766=>x"000c5",
2767=>x"000c5",
2768=>x"000c5",
2769=>x"000c5",
2770=>x"000c5",
2771=>x"000c5",
2772=>x"000c6",
2773=>x"000c6",
2774=>x"000c6",
2775=>x"000c6",
2776=>x"000c6",
2777=>x"000c6",
2778=>x"000c6",
2779=>x"000c6",
2780=>x"000c6",
2781=>x"000c6",
2782=>x"000c6",
2783=>x"000c6",
2784=>x"000c6",
2785=>x"000c6",
2786=>x"000c7",
2787=>x"000c7",
2788=>x"000c7",
2789=>x"000c7",
2790=>x"000c7",
2791=>x"000c7",
2792=>x"000c7",
2793=>x"000c7",
2794=>x"000c7",
2795=>x"000c7",
2796=>x"000c7",
2797=>x"000c7",
2798=>x"000c7",
2799=>x"000c7",
2800=>x"000c8",
2801=>x"000c8",
2802=>x"000c8",
2803=>x"000c8",
2804=>x"000c8",
2805=>x"000c8",
2806=>x"000c8",
2807=>x"000c8",
2808=>x"000c8",
2809=>x"000c8",
2810=>x"000c8",
2811=>x"000c8",
2812=>x"000c8",
2813=>x"000c8",
2814=>x"000c9",
2815=>x"000c9",
2816=>x"000c9",
2817=>x"000c9",
2818=>x"000c9",
2819=>x"000c9",
2820=>x"000c9",
2821=>x"000c9",
2822=>x"000c9",
2823=>x"000c9",
2824=>x"000c9",
2825=>x"000c9",
2826=>x"000c9",
2827=>x"000c9",
2828=>x"000ca",
2829=>x"000ca",
2830=>x"000ca",
2831=>x"000ca",
2832=>x"000ca",
2833=>x"000ca",
2834=>x"000ca",
2835=>x"000ca",
2836=>x"000ca",
2837=>x"000ca",
2838=>x"000ca",
2839=>x"000ca",
2840=>x"000ca",
2841=>x"000ca",
2842=>x"000cb",
2843=>x"000cb",
2844=>x"000cb",
2845=>x"000cb",
2846=>x"000cb",
2847=>x"000cb",
2848=>x"000cb",
2849=>x"000cb",
2850=>x"000cb",
2851=>x"000cb",
2852=>x"000cb",
2853=>x"000cb",
2854=>x"000cb",
2855=>x"000cb",
2856=>x"000cc",
2857=>x"000cc",
2858=>x"000cc",
2859=>x"000cc",
2860=>x"000cc",
2861=>x"000cc",
2862=>x"000cc",
2863=>x"000cc",
2864=>x"000cc",
2865=>x"000cc",
2866=>x"000cc",
2867=>x"000cc",
2868=>x"000cc",
2869=>x"000cc",
2870=>x"000cd",
2871=>x"000cd",
2872=>x"000cd",
2873=>x"000cd",
2874=>x"000cd",
2875=>x"000cd",
2876=>x"000cd",
2877=>x"000cd",
2878=>x"000cd",
2879=>x"000cd",
2880=>x"000cd",
2881=>x"000cd",
2882=>x"000cd",
2883=>x"000cd",
2884=>x"000ce",
2885=>x"000ce",
2886=>x"000ce",
2887=>x"000ce",
2888=>x"000ce",
2889=>x"000ce",
2890=>x"000ce",
2891=>x"000ce",
2892=>x"000ce",
2893=>x"000ce",
2894=>x"000ce",
2895=>x"000ce",
2896=>x"000ce",
2897=>x"000ce",
2898=>x"000cf",
2899=>x"000cf",
2900=>x"000cf",
2901=>x"000cf",
2902=>x"000cf",
2903=>x"000cf",
2904=>x"000cf",
2905=>x"000cf",
2906=>x"000cf",
2907=>x"000cf",
2908=>x"000cf",
2909=>x"000cf",
2910=>x"000cf",
2911=>x"000cf",
2912=>x"000d0",
2913=>x"000d0",
2914=>x"000d0",
2915=>x"000d0",
2916=>x"000d0",
2917=>x"000d0",
2918=>x"000d0",
2919=>x"000d0",
2920=>x"000d0",
2921=>x"000d0",
2922=>x"000d0",
2923=>x"000d0",
2924=>x"000d0",
2925=>x"000d0",
2926=>x"000d1",
2927=>x"000d1",
2928=>x"000d1",
2929=>x"000d1",
2930=>x"000d1",
2931=>x"000d1",
2932=>x"000d1",
2933=>x"000d1",
2934=>x"000d1",
2935=>x"000d1",
2936=>x"000d1",
2937=>x"000d1",
2938=>x"000d1",
2939=>x"000d1",
2940=>x"000d2",
2941=>x"000d2",
2942=>x"000d2",
2943=>x"000d2",
2944=>x"000d2",
2945=>x"000d2",
2946=>x"000d2",
2947=>x"000d2",
2948=>x"000d2",
2949=>x"000d2",
2950=>x"000d2",
2951=>x"000d2",
2952=>x"000d2",
2953=>x"000d2",
2954=>x"000d3",
2955=>x"000d3",
2956=>x"000d3",
2957=>x"000d3",
2958=>x"000d3",
2959=>x"000d3",
2960=>x"000d3",
2961=>x"000d3",
2962=>x"000d3",
2963=>x"000d3",
2964=>x"000d3",
2965=>x"000d3",
2966=>x"000d3",
2967=>x"000d3",
2968=>x"000d4",
2969=>x"000d4",
2970=>x"000d4",
2971=>x"000d4",
2972=>x"000d4",
2973=>x"000d4",
2974=>x"000d4",
2975=>x"000d4",
2976=>x"000d4",
2977=>x"000d4",
2978=>x"000d4",
2979=>x"000d4",
2980=>x"000d4",
2981=>x"000d4",
2982=>x"000d5",
2983=>x"000d5",
2984=>x"000d5",
2985=>x"000d5",
2986=>x"000d5",
2987=>x"000d5",
2988=>x"000d5",
2989=>x"000d5",
2990=>x"000d5",
2991=>x"000d5",
2992=>x"000d5",
2993=>x"000d5",
2994=>x"000d5",
2995=>x"000d5",
2996=>x"000d6",
2997=>x"000d6",
2998=>x"000d6",
2999=>x"000d6",
3000=>x"000d6",
3001=>x"000d6",
3002=>x"000d6",
3003=>x"000d6",
3004=>x"000d6",
3005=>x"000d6",
3006=>x"000d6",
3007=>x"000d6",
3008=>x"000d6",
3009=>x"000d6",
3010=>x"000d7",
3011=>x"000d7",
3012=>x"000d7",
3013=>x"000d7",
3014=>x"000d7",
3015=>x"000d7",
3016=>x"000d7",
3017=>x"000d7",
3018=>x"000d7",
3019=>x"000d7",
3020=>x"000d7",
3021=>x"000d7",
3022=>x"000d7",
3023=>x"000d7",
3024=>x"000d8",
3025=>x"000d8",
3026=>x"000d8",
3027=>x"000d8",
3028=>x"000d8",
3029=>x"000d8",
3030=>x"000d8",
3031=>x"000d8",
3032=>x"000d8",
3033=>x"000d8",
3034=>x"000d8",
3035=>x"000d8",
3036=>x"000d8",
3037=>x"000d8",
3038=>x"000d9",
3039=>x"000d9",
3040=>x"000d9",
3041=>x"000d9",
3042=>x"000d9",
3043=>x"000d9",
3044=>x"000d9",
3045=>x"000d9",
3046=>x"000d9",
3047=>x"000d9",
3048=>x"000d9",
3049=>x"000d9",
3050=>x"000d9",
3051=>x"000d9",
3052=>x"000da",
3053=>x"000da",
3054=>x"000da",
3055=>x"000da",
3056=>x"000da",
3057=>x"000da",
3058=>x"000da",
3059=>x"000da",
3060=>x"000da",
3061=>x"000da",
3062=>x"000da",
3063=>x"000da",
3064=>x"000da",
3065=>x"000da",
3066=>x"000db",
3067=>x"000db",
3068=>x"000db",
3069=>x"000db",
3070=>x"000db",
3071=>x"000db",
3072=>x"000db",
3073=>x"000db",
3074=>x"000db",
3075=>x"000db",
3076=>x"000db",
3077=>x"000db",
3078=>x"000db",
3079=>x"000db",
3080=>x"000dc",
3081=>x"000dc",
3082=>x"000dc",
3083=>x"000dc",
3084=>x"000dc",
3085=>x"000dc",
3086=>x"000dc",
3087=>x"000dc",
3088=>x"000dc",
3089=>x"000dc",
3090=>x"000dc",
3091=>x"000dc",
3092=>x"000dc",
3093=>x"000dc",
3094=>x"000dd",
3095=>x"000dd",
3096=>x"000dd",
3097=>x"000dd",
3098=>x"000dd",
3099=>x"000dd",
3100=>x"000dd",
3101=>x"000dd",
3102=>x"000dd",
3103=>x"000dd",
3104=>x"000dd",
3105=>x"000dd",
3106=>x"000dd",
3107=>x"000dd",
3108=>x"000de",
3109=>x"000de",
3110=>x"000de",
3111=>x"000de",
3112=>x"000de",
3113=>x"000de",
3114=>x"000de",
3115=>x"000de",
3116=>x"000de",
3117=>x"000de",
3118=>x"000de",
3119=>x"000de",
3120=>x"000de",
3121=>x"000de",
3122=>x"000df",
3123=>x"000df",
3124=>x"000df",
3125=>x"000df",
3126=>x"000df",
3127=>x"000df",
3128=>x"000df",
3129=>x"000df",
3130=>x"000df",
3131=>x"000df",
3132=>x"000df",
3133=>x"000df",
3134=>x"000df",
3135=>x"000df",
3136=>x"000e0",
3137=>x"000e0",
3138=>x"000e0",
3139=>x"000e0",
3140=>x"000e0",
3141=>x"000e0",
3142=>x"000e0",
3143=>x"000e0",
3144=>x"000e0",
3145=>x"000e0",
3146=>x"000e0",
3147=>x"000e0",
3148=>x"000e0",
3149=>x"000e0",
3150=>x"000e1",
3151=>x"000e1",
3152=>x"000e1",
3153=>x"000e1",
3154=>x"000e1",
3155=>x"000e1",
3156=>x"000e1",
3157=>x"000e1",
3158=>x"000e1",
3159=>x"000e1",
3160=>x"000e1",
3161=>x"000e1",
3162=>x"000e1",
3163=>x"000e1",
3164=>x"000e2",
3165=>x"000e2",
3166=>x"000e2",
3167=>x"000e2",
3168=>x"000e2",
3169=>x"000e2",
3170=>x"000e2",
3171=>x"000e2",
3172=>x"000e2",
3173=>x"000e2",
3174=>x"000e2",
3175=>x"000e2",
3176=>x"000e2",
3177=>x"000e2",
3178=>x"000e3",
3179=>x"000e3",
3180=>x"000e3",
3181=>x"000e3",
3182=>x"000e3",
3183=>x"000e3",
3184=>x"000e3",
3185=>x"000e3",
3186=>x"000e3",
3187=>x"000e3",
3188=>x"000e3",
3189=>x"000e3",
3190=>x"000e3",
3191=>x"000e3",
3192=>x"000e4",
3193=>x"000e4",
3194=>x"000e4",
3195=>x"000e4",
3196=>x"000e4",
3197=>x"000e4",
3198=>x"000e4",
3199=>x"000e4",
3200=>x"000e4",
3201=>x"000e4",
3202=>x"000e4",
3203=>x"000e4",
3204=>x"000e4",
3205=>x"000e4",
3206=>x"000e5",
3207=>x"000e5",
3208=>x"000e5",
3209=>x"000e5",
3210=>x"000e5",
3211=>x"000e5",
3212=>x"000e5",
3213=>x"000e5",
3214=>x"000e5",
3215=>x"000e5",
3216=>x"000e5",
3217=>x"000e5",
3218=>x"000e5",
3219=>x"000e5",
3220=>x"000e6",
3221=>x"000e6",
3222=>x"000e6",
3223=>x"000e6",
3224=>x"000e6",
3225=>x"000e6",
3226=>x"000e6",
3227=>x"000e6",
3228=>x"000e6",
3229=>x"000e6",
3230=>x"000e6",
3231=>x"000e6",
3232=>x"000e6",
3233=>x"000e6",
3234=>x"000e7",
3235=>x"000e7",
3236=>x"000e7",
3237=>x"000e7",
3238=>x"000e7",
3239=>x"000e7",
3240=>x"000e7",
3241=>x"000e7",
3242=>x"000e7",
3243=>x"000e7",
3244=>x"000e7",
3245=>x"000e7",
3246=>x"000e7",
3247=>x"000e7",
3248=>x"000e8",
3249=>x"000e8",
3250=>x"000e8",
3251=>x"000e8",
3252=>x"000e8",
3253=>x"000e8",
3254=>x"000e8",
3255=>x"000e8",
3256=>x"000e8",
3257=>x"000e8",
3258=>x"000e8",
3259=>x"000e8",
3260=>x"000e8",
3261=>x"000e8",
3262=>x"000e9",
3263=>x"000e9",
3264=>x"000e9",
3265=>x"000e9",
3266=>x"000e9",
3267=>x"000e9",
3268=>x"000e9",
3269=>x"000e9",
3270=>x"000e9",
3271=>x"000e9",
3272=>x"000e9",
3273=>x"000e9",
3274=>x"000e9",
3275=>x"000e9",
3276=>x"000ea",
3277=>x"000ea",
3278=>x"000ea",
3279=>x"000ea",
3280=>x"000ea",
3281=>x"000ea",
3282=>x"000ea",
3283=>x"000ea",
3284=>x"000ea",
3285=>x"000ea",
3286=>x"000ea",
3287=>x"000ea",
3288=>x"000ea",
3289=>x"000ea",
3290=>x"000eb",
3291=>x"000eb",
3292=>x"000eb",
3293=>x"000eb",
3294=>x"000eb",
3295=>x"000eb",
3296=>x"000eb",
3297=>x"000eb",
3298=>x"000eb",
3299=>x"000eb",
3300=>x"000eb",
3301=>x"000eb",
3302=>x"000eb",
3303=>x"000eb",
3304=>x"000ec",
3305=>x"000ec",
3306=>x"000ec",
3307=>x"000ec",
3308=>x"000ec",
3309=>x"000ec",
3310=>x"000ec",
3311=>x"000ec",
3312=>x"000ec",
3313=>x"000ec",
3314=>x"000ec",
3315=>x"000ec",
3316=>x"000ec",
3317=>x"000ec",
3318=>x"000ed",
3319=>x"000ed",
3320=>x"000ed",
3321=>x"000ed",
3322=>x"000ed",
3323=>x"000ed",
3324=>x"000ed",
3325=>x"000ed",
3326=>x"000ed",
3327=>x"000ed",
3328=>x"000ed",
3329=>x"000ed",
3330=>x"000ed",
3331=>x"000ed",
3332=>x"000ee",
3333=>x"000ee",
3334=>x"000ee",
3335=>x"000ee",
3336=>x"000ee",
3337=>x"000ee",
3338=>x"000ee",
3339=>x"000ee",
3340=>x"000ee",
3341=>x"000ee",
3342=>x"000ee",
3343=>x"000ee",
3344=>x"000ee",
3345=>x"000ee",
3346=>x"000ef",
3347=>x"000ef",
3348=>x"000ef",
3349=>x"000ef",
3350=>x"000ef",
3351=>x"000ef",
3352=>x"000ef",
3353=>x"000ef",
3354=>x"000ef",
3355=>x"000ef",
3356=>x"000ef",
3357=>x"000ef",
3358=>x"000ef",
3359=>x"000ef",
3360=>x"000f0",
3361=>x"000f0",
3362=>x"000f0",
3363=>x"000f0",
3364=>x"000f0",
3365=>x"000f0",
3366=>x"000f0",
3367=>x"000f0",
3368=>x"000f0",
3369=>x"000f0",
3370=>x"000f0",
3371=>x"000f0",
3372=>x"000f0",
3373=>x"000f0",
3374=>x"000f1",
3375=>x"000f1",
3376=>x"000f1",
3377=>x"000f1",
3378=>x"000f1",
3379=>x"000f1",
3380=>x"000f1",
3381=>x"000f1",
3382=>x"000f1",
3383=>x"000f1",
3384=>x"000f1",
3385=>x"000f1",
3386=>x"000f1",
3387=>x"000f1",
3388=>x"000f2",
3389=>x"000f2",
3390=>x"000f2",
3391=>x"000f2",
3392=>x"000f2",
3393=>x"000f2",
3394=>x"000f2",
3395=>x"000f2",
3396=>x"000f2",
3397=>x"000f2",
3398=>x"000f2",
3399=>x"000f2",
3400=>x"000f2",
3401=>x"000f2",
3402=>x"000f3",
3403=>x"000f3",
3404=>x"000f3",
3405=>x"000f3",
3406=>x"000f3",
3407=>x"000f3",
3408=>x"000f3",
3409=>x"000f3",
3410=>x"000f3",
3411=>x"000f3",
3412=>x"000f3",
3413=>x"000f3",
3414=>x"000f3",
3415=>x"000f3",
3416=>x"000f4",
3417=>x"000f4",
3418=>x"000f4",
3419=>x"000f4",
3420=>x"000f4",
3421=>x"000f4",
3422=>x"000f4",
3423=>x"000f4",
3424=>x"000f4",
3425=>x"000f4",
3426=>x"000f4",
3427=>x"000f4",
3428=>x"000f4",
3429=>x"000f4",
3430=>x"000f5",
3431=>x"000f5",
3432=>x"000f5",
3433=>x"000f5",
3434=>x"000f5",
3435=>x"000f5",
3436=>x"000f5",
3437=>x"000f5",
3438=>x"000f5",
3439=>x"000f5",
3440=>x"000f5",
3441=>x"000f5",
3442=>x"000f5",
3443=>x"000f5",
3444=>x"000f6",
3445=>x"000f6",
3446=>x"000f6",
3447=>x"000f6",
3448=>x"000f6",
3449=>x"000f6",
3450=>x"000f6",
3451=>x"000f6",
3452=>x"000f6",
3453=>x"000f6",
3454=>x"000f6",
3455=>x"000f6",
3456=>x"000f6",
3457=>x"000f6",
3458=>x"000f7",
3459=>x"000f7",
3460=>x"000f7",
3461=>x"000f7",
3462=>x"000f7",
3463=>x"000f7",
3464=>x"000f7",
3465=>x"000f7",
3466=>x"000f7",
3467=>x"000f7",
3468=>x"000f7",
3469=>x"000f7",
3470=>x"000f7",
3471=>x"000f7",
3472=>x"000f8",
3473=>x"000f8",
3474=>x"000f8",
3475=>x"000f8",
3476=>x"000f8",
3477=>x"000f8",
3478=>x"000f8",
3479=>x"000f8",
3480=>x"000f8",
3481=>x"000f8",
3482=>x"000f8",
3483=>x"000f8",
3484=>x"000f8",
3485=>x"000f8",
3486=>x"000f9",
3487=>x"000f9",
3488=>x"000f9",
3489=>x"000f9",
3490=>x"000f9",
3491=>x"000f9",
3492=>x"000f9",
3493=>x"000f9",
3494=>x"000f9",
3495=>x"000f9",
3496=>x"000f9",
3497=>x"000f9",
3498=>x"000f9",
3499=>x"000f9",
3500=>x"000fa",
3501=>x"000fa",
3502=>x"000fa",
3503=>x"000fa",
3504=>x"000fa",
3505=>x"000fa",
3506=>x"000fa",
3507=>x"000fa",
3508=>x"000fa",
3509=>x"000fa",
3510=>x"000fa",
3511=>x"000fa",
3512=>x"000fa",
3513=>x"000fa",
3514=>x"000fb",
3515=>x"000fb",
3516=>x"000fb",
3517=>x"000fb",
3518=>x"000fb",
3519=>x"000fb",
3520=>x"000fb",
3521=>x"000fb",
3522=>x"000fb",
3523=>x"000fb",
3524=>x"000fb",
3525=>x"000fb",
3526=>x"000fb",
3527=>x"000fb",
3528=>x"000fc",
3529=>x"000fc",
3530=>x"000fc",
3531=>x"000fc",
3532=>x"000fc",
3533=>x"000fc",
3534=>x"000fc",
3535=>x"000fc",
3536=>x"000fc",
3537=>x"000fc",
3538=>x"000fc",
3539=>x"000fc",
3540=>x"000fc",
3541=>x"000fc",
3542=>x"000fd",
3543=>x"000fd",
3544=>x"000fd",
3545=>x"000fd",
3546=>x"000fd",
3547=>x"000fd",
3548=>x"000fd",
3549=>x"000fd",
3550=>x"000fd",
3551=>x"000fd",
3552=>x"000fd",
3553=>x"000fd",
3554=>x"000fd",
3555=>x"000fd",
3556=>x"000fe",
3557=>x"000fe",
3558=>x"000fe",
3559=>x"000fe",
3560=>x"000fe",
3561=>x"000fe",
3562=>x"000fe",
3563=>x"000fe",
3564=>x"000fe",
3565=>x"000fe",
3566=>x"000fe",
3567=>x"000fe",
3568=>x"000fe",
3569=>x"000fe",
3570=>x"000ff",
3571=>x"000ff",
3572=>x"000ff",
3573=>x"000ff",
3574=>x"000ff",
3575=>x"000ff",
3576=>x"000ff",
3577=>x"000ff",
3578=>x"000ff",
3579=>x"000ff",
3580=>x"000ff",
3581=>x"000ff",
3582=>x"000ff",
3583=>x"000ff",
3584=>x"00100",
3585=>x"00100",
3586=>x"00100",
3587=>x"00100",
3588=>x"00100",
3589=>x"00100",
3590=>x"00100",
3591=>x"00100",
3592=>x"00100",
3593=>x"00100",
3594=>x"00100",
3595=>x"00100",
3596=>x"00100",
3597=>x"00100",
3598=>x"00101",
3599=>x"00101",
3600=>x"00101",
3601=>x"00101",
3602=>x"00101",
3603=>x"00101",
3604=>x"00101",
3605=>x"00101",
3606=>x"00101",
3607=>x"00101",
3608=>x"00101",
3609=>x"00101",
3610=>x"00101",
3611=>x"00101",
3612=>x"00102",
3613=>x"00102",
3614=>x"00102",
3615=>x"00102",
3616=>x"00102",
3617=>x"00102",
3618=>x"00102",
3619=>x"00102",
3620=>x"00102",
3621=>x"00102",
3622=>x"00102",
3623=>x"00102",
3624=>x"00102",
3625=>x"00102",
3626=>x"00103",
3627=>x"00103",
3628=>x"00103",
3629=>x"00103",
3630=>x"00103",
3631=>x"00103",
3632=>x"00103",
3633=>x"00103",
3634=>x"00103",
3635=>x"00103",
3636=>x"00103",
3637=>x"00103",
3638=>x"00103",
3639=>x"00103",
3640=>x"00104",
3641=>x"00104",
3642=>x"00104",
3643=>x"00104",
3644=>x"00104",
3645=>x"00104",
3646=>x"00104",
3647=>x"00104",
3648=>x"00104",
3649=>x"00104",
3650=>x"00104",
3651=>x"00104",
3652=>x"00104",
3653=>x"00104",
3654=>x"00105",
3655=>x"00105",
3656=>x"00105",
3657=>x"00105",
3658=>x"00105",
3659=>x"00105",
3660=>x"00105",
3661=>x"00105",
3662=>x"00105",
3663=>x"00105",
3664=>x"00105",
3665=>x"00105",
3666=>x"00105",
3667=>x"00105",
3668=>x"00106",
3669=>x"00106",
3670=>x"00106",
3671=>x"00106",
3672=>x"00106",
3673=>x"00106",
3674=>x"00106",
3675=>x"00106",
3676=>x"00106",
3677=>x"00106",
3678=>x"00106",
3679=>x"00106",
3680=>x"00106",
3681=>x"00106",
3682=>x"00107",
3683=>x"00107",
3684=>x"00107",
3685=>x"00107",
3686=>x"00107",
3687=>x"00107",
3688=>x"00107",
3689=>x"00107",
3690=>x"00107",
3691=>x"00107",
3692=>x"00107",
3693=>x"00107",
3694=>x"00107",
3695=>x"00107",
3696=>x"00108",
3697=>x"00108",
3698=>x"00108",
3699=>x"00108",
3700=>x"00108",
3701=>x"00108",
3702=>x"00108",
3703=>x"00108",
3704=>x"00108",
3705=>x"00108",
3706=>x"00108",
3707=>x"00108",
3708=>x"00108",
3709=>x"00108",
3710=>x"00109",
3711=>x"00109",
3712=>x"00109",
3713=>x"00109",
3714=>x"00109",
3715=>x"00109",
3716=>x"00109",
3717=>x"00109",
3718=>x"00109",
3719=>x"00109",
3720=>x"00109",
3721=>x"00109",
3722=>x"00109",
3723=>x"00109",
3724=>x"0010a",
3725=>x"0010a",
3726=>x"0010a",
3727=>x"0010a",
3728=>x"0010a",
3729=>x"0010a",
3730=>x"0010a",
3731=>x"0010a",
3732=>x"0010a",
3733=>x"0010a",
3734=>x"0010a",
3735=>x"0010a",
3736=>x"0010a",
3737=>x"0010a",
3738=>x"0010b",
3739=>x"0010b",
3740=>x"0010b",
3741=>x"0010b",
3742=>x"0010b",
3743=>x"0010b",
3744=>x"0010b",
3745=>x"0010b",
3746=>x"0010b",
3747=>x"0010b",
3748=>x"0010b",
3749=>x"0010b",
3750=>x"0010b",
3751=>x"0010b",
3752=>x"0010c",
3753=>x"0010c",
3754=>x"0010c",
3755=>x"0010c",
3756=>x"0010c",
3757=>x"0010c",
3758=>x"0010c",
3759=>x"0010c",
3760=>x"0010c",
3761=>x"0010c",
3762=>x"0010c",
3763=>x"0010c",
3764=>x"0010c",
3765=>x"0010c",
3766=>x"0010d",
3767=>x"0010d",
3768=>x"0010d",
3769=>x"0010d",
3770=>x"0010d",
3771=>x"0010d",
3772=>x"0010d",
3773=>x"0010d",
3774=>x"0010d",
3775=>x"0010d",
3776=>x"0010d",
3777=>x"0010d",
3778=>x"0010d",
3779=>x"0010d",
3780=>x"0010e",
3781=>x"0010e",
3782=>x"0010e",
3783=>x"0010e",
3784=>x"0010e",
3785=>x"0010e",
3786=>x"0010e",
3787=>x"0010e",
3788=>x"0010e",
3789=>x"0010e",
3790=>x"0010e",
3791=>x"0010e",
3792=>x"0010e",
3793=>x"0010e",
3794=>x"0010f",
3795=>x"0010f",
3796=>x"0010f",
3797=>x"0010f",
3798=>x"0010f",
3799=>x"0010f",
3800=>x"0010f",
3801=>x"0010f",
3802=>x"0010f",
3803=>x"0010f",
3804=>x"0010f",
3805=>x"0010f",
3806=>x"0010f",
3807=>x"0010f",
3808=>x"00110",
3809=>x"00110",
3810=>x"00110",
3811=>x"00110",
3812=>x"00110",
3813=>x"00110",
3814=>x"00110",
3815=>x"00110",
3816=>x"00110",
3817=>x"00110",
3818=>x"00110",
3819=>x"00110",
3820=>x"00110",
3821=>x"00110",
3822=>x"00111",
3823=>x"00111",
3824=>x"00111",
3825=>x"00111",
3826=>x"00111",
3827=>x"00111",
3828=>x"00111",
3829=>x"00111",
3830=>x"00111",
3831=>x"00111",
3832=>x"00111",
3833=>x"00111",
3834=>x"00111",
3835=>x"00111",
3836=>x"00112",
3837=>x"00112",
3838=>x"00112",
3839=>x"00112",
3840=>x"00112",
3841=>x"00112",
3842=>x"00112",
3843=>x"00112",
3844=>x"00112",
3845=>x"00112",
3846=>x"00112",
3847=>x"00112",
3848=>x"00112",
3849=>x"00112",
3850=>x"00113",
3851=>x"00113",
3852=>x"00113",
3853=>x"00113",
3854=>x"00113",
3855=>x"00113",
3856=>x"00113",
3857=>x"00113",
3858=>x"00113",
3859=>x"00113",
3860=>x"00113",
3861=>x"00113",
3862=>x"00113",
3863=>x"00113",
3864=>x"00114",
3865=>x"00114",
3866=>x"00114",
3867=>x"00114",
3868=>x"00114",
3869=>x"00114",
3870=>x"00114",
3871=>x"00114",
3872=>x"00114",
3873=>x"00114",
3874=>x"00114",
3875=>x"00114",
3876=>x"00114",
3877=>x"00114",
3878=>x"00115",
3879=>x"00115",
3880=>x"00115",
3881=>x"00115",
3882=>x"00115",
3883=>x"00115",
3884=>x"00115",
3885=>x"00115",
3886=>x"00115",
3887=>x"00115",
3888=>x"00115",
3889=>x"00115",
3890=>x"00115",
3891=>x"00115",
3892=>x"00116",
3893=>x"00116",
3894=>x"00116",
3895=>x"00116",
3896=>x"00116",
3897=>x"00116",
3898=>x"00116",
3899=>x"00116",
3900=>x"00116",
3901=>x"00116",
3902=>x"00116",
3903=>x"00116",
3904=>x"00116",
3905=>x"00116",
3906=>x"00117",
3907=>x"00117",
3908=>x"00117",
3909=>x"00117",
3910=>x"00117",
3911=>x"00117",
3912=>x"00117",
3913=>x"00117",
3914=>x"00117",
3915=>x"00117",
3916=>x"00117",
3917=>x"00117",
3918=>x"00117",
3919=>x"00117",
3920=>x"00118",
3921=>x"00118",
3922=>x"00118",
3923=>x"00118",
3924=>x"00118",
3925=>x"00118",
3926=>x"00118",
3927=>x"00118",
3928=>x"00118",
3929=>x"00118",
3930=>x"00118",
3931=>x"00118",
3932=>x"00118",
3933=>x"00118",
3934=>x"00119",
3935=>x"00119",
3936=>x"00119",
3937=>x"00119",
3938=>x"00119",
3939=>x"00119",
3940=>x"00119",
3941=>x"00119",
3942=>x"00119",
3943=>x"00119",
3944=>x"00119",
3945=>x"00119",
3946=>x"00119",
3947=>x"00119",
3948=>x"0011a",
3949=>x"0011a",
3950=>x"0011a",
3951=>x"0011a",
3952=>x"0011a",
3953=>x"0011a",
3954=>x"0011a",
3955=>x"0011a",
3956=>x"0011a",
3957=>x"0011a",
3958=>x"0011a",
3959=>x"0011a",
3960=>x"0011a",
3961=>x"0011a",
3962=>x"0011b",
3963=>x"0011b",
3964=>x"0011b",
3965=>x"0011b",
3966=>x"0011b",
3967=>x"0011b",
3968=>x"0011b",
3969=>x"0011b",
3970=>x"0011b",
3971=>x"0011b",
3972=>x"0011b",
3973=>x"0011b",
3974=>x"0011b",
3975=>x"0011b",
3976=>x"0011c",
3977=>x"0011c",
3978=>x"0011c",
3979=>x"0011c",
3980=>x"0011c",
3981=>x"0011c",
3982=>x"0011c",
3983=>x"0011c",
3984=>x"0011c",
3985=>x"0011c",
3986=>x"0011c",
3987=>x"0011c",
3988=>x"0011c",
3989=>x"0011c",
3990=>x"0011d",
3991=>x"0011d",
3992=>x"0011d",
3993=>x"0011d",
3994=>x"0011d",
3995=>x"0011d",
3996=>x"0011d",
3997=>x"0011d",
3998=>x"0011d",
3999=>x"0011d",
4000=>x"0011d",
4001=>x"0011d",
4002=>x"0011d",
4003=>x"0011d",
4004=>x"0011e",
4005=>x"0011e",
4006=>x"0011e",
4007=>x"0011e",
4008=>x"0011e",
4009=>x"0011e",
4010=>x"0011e",
4011=>x"0011e",
4012=>x"0011e",
4013=>x"0011e",
4014=>x"0011e",
4015=>x"0011e",
4016=>x"0011e",
4017=>x"0011e",
4018=>x"0011f",
4019=>x"0011f",
4020=>x"0011f",
4021=>x"0011f",
4022=>x"0011f",
4023=>x"0011f",
4024=>x"0011f",
4025=>x"0011f",
4026=>x"0011f",
4027=>x"0011f",
4028=>x"0011f",
4029=>x"0011f",
4030=>x"0011f",
4031=>x"0011f",
4032=>x"00120",
4033=>x"00120",
4034=>x"00120",
4035=>x"00120",
4036=>x"00120",
4037=>x"00120",
4038=>x"00120",
4039=>x"00120",
4040=>x"00120",
4041=>x"00120",
4042=>x"00120",
4043=>x"00120",
4044=>x"00120",
4045=>x"00120",
4046=>x"00121",
4047=>x"00121",
4048=>x"00121",
4049=>x"00121",
4050=>x"00121",
4051=>x"00121",
4052=>x"00121",
4053=>x"00121",
4054=>x"00121",
4055=>x"00121",
4056=>x"00121",
4057=>x"00121",
4058=>x"00121",
4059=>x"00121",
4060=>x"00122",
4061=>x"00122",
4062=>x"00122",
4063=>x"00122",
4064=>x"00122",
4065=>x"00122",
4066=>x"00122",
4067=>x"00122",
4068=>x"00122",
4069=>x"00122",
4070=>x"00122",
4071=>x"00122",
4072=>x"00122",
4073=>x"00122",
4074=>x"00123",
4075=>x"00123",
4076=>x"00123",
4077=>x"00123",
4078=>x"00123",
4079=>x"00123",
4080=>x"00123",
4081=>x"00123",
4082=>x"00123",
4083=>x"00123",
4084=>x"00123",
4085=>x"00123",
4086=>x"00123",
4087=>x"00123",
4088=>x"00124",
4089=>x"00124",
4090=>x"00124",
4091=>x"00124",
4092=>x"00124",
4093=>x"00124",
4094=>x"00124",
4095=>x"00124",
4096=>x"00124",
4097=>x"00124",
4098=>x"00124",
4099=>x"00124",
4100=>x"00124",
4101=>x"00124",
4102=>x"00125",
4103=>x"00125",
4104=>x"00125",
4105=>x"00125",
4106=>x"00125",
4107=>x"00125",
4108=>x"00125",
4109=>x"00125",
4110=>x"00125",
4111=>x"00125",
4112=>x"00125",
4113=>x"00125",
4114=>x"00125",
4115=>x"00125",
4116=>x"00126",
4117=>x"00126",
4118=>x"00126",
4119=>x"00126",
4120=>x"00126",
4121=>x"00126",
4122=>x"00126",
4123=>x"00126",
4124=>x"00126",
4125=>x"00126",
4126=>x"00126",
4127=>x"00126",
4128=>x"00126",
4129=>x"00126",
4130=>x"00127",
4131=>x"00127",
4132=>x"00127",
4133=>x"00127",
4134=>x"00127",
4135=>x"00127",
4136=>x"00127",
4137=>x"00127",
4138=>x"00127",
4139=>x"00127",
4140=>x"00127",
4141=>x"00127",
4142=>x"00127",
4143=>x"00127",
4144=>x"00128",
4145=>x"00128",
4146=>x"00128",
4147=>x"00128",
4148=>x"00128",
4149=>x"00128",
4150=>x"00128",
4151=>x"00128",
4152=>x"00128",
4153=>x"00128",
4154=>x"00128",
4155=>x"00128",
4156=>x"00128",
4157=>x"00128",
4158=>x"00129",
4159=>x"00129",
4160=>x"00129",
4161=>x"00129",
4162=>x"00129",
4163=>x"00129",
4164=>x"00129",
4165=>x"00129",
4166=>x"00129",
4167=>x"00129",
4168=>x"00129",
4169=>x"00129",
4170=>x"00129",
4171=>x"00129",
4172=>x"0012a",
4173=>x"0012a",
4174=>x"0012a",
4175=>x"0012a",
4176=>x"0012a",
4177=>x"0012a",
4178=>x"0012a",
4179=>x"0012a",
4180=>x"0012a",
4181=>x"0012a",
4182=>x"0012a",
4183=>x"0012a",
4184=>x"0012a",
4185=>x"0012a",
4186=>x"0012b",
4187=>x"0012b",
4188=>x"0012b",
4189=>x"0012b",
4190=>x"0012b",
4191=>x"0012b",
4192=>x"0012b",
4193=>x"0012b",
4194=>x"0012b",
4195=>x"0012b",
4196=>x"0012b",
4197=>x"0012b",
4198=>x"0012b",
4199=>x"0012b",
4200=>x"0012c",
4201=>x"0012c",
4202=>x"0012c",
4203=>x"0012c",
4204=>x"0012c",
4205=>x"0012c",
4206=>x"0012c",
4207=>x"0012c",
4208=>x"0012c",
4209=>x"0012c",
4210=>x"0012c",
4211=>x"0012c",
4212=>x"0012c",
4213=>x"0012c",
4214=>x"0012d",
4215=>x"0012d",
4216=>x"0012d",
4217=>x"0012d",
4218=>x"0012d",
4219=>x"0012d",
4220=>x"0012d",
4221=>x"0012d",
4222=>x"0012d",
4223=>x"0012d",
4224=>x"0012d",
4225=>x"0012d",
4226=>x"0012d",
4227=>x"0012d",
4228=>x"0012e",
4229=>x"0012e",
4230=>x"0012e",
4231=>x"0012e",
4232=>x"0012e",
4233=>x"0012e",
4234=>x"0012e",
4235=>x"0012e",
4236=>x"0012e",
4237=>x"0012e",
4238=>x"0012e",
4239=>x"0012e",
4240=>x"0012e",
4241=>x"0012e",
4242=>x"0012f",
4243=>x"0012f",
4244=>x"0012f",
4245=>x"0012f",
4246=>x"0012f",
4247=>x"0012f",
4248=>x"0012f",
4249=>x"0012f",
4250=>x"0012f",
4251=>x"0012f",
4252=>x"0012f",
4253=>x"0012f",
4254=>x"0012f",
4255=>x"0012f",
4256=>x"00130",
4257=>x"00130",
4258=>x"00130",
4259=>x"00130",
4260=>x"00130",
4261=>x"00130",
4262=>x"00130",
4263=>x"00130",
4264=>x"00130",
4265=>x"00130",
4266=>x"00130",
4267=>x"00130",
4268=>x"00130",
4269=>x"00130",
4270=>x"00131",
4271=>x"00131",
4272=>x"00131",
4273=>x"00131",
4274=>x"00131",
4275=>x"00131",
4276=>x"00131",
4277=>x"00131",
4278=>x"00131",
4279=>x"00131",
4280=>x"00131",
4281=>x"00131",
4282=>x"00131",
4283=>x"00131",
4284=>x"00132",
4285=>x"00132",
4286=>x"00132",
4287=>x"00132",
4288=>x"00132",
4289=>x"00132",
4290=>x"00132",
4291=>x"00132",
4292=>x"00132",
4293=>x"00132",
4294=>x"00132",
4295=>x"00132",
4296=>x"00132",
4297=>x"00132",
4298=>x"00133",
4299=>x"00133",
4300=>x"00133",
4301=>x"00133",
4302=>x"00133",
4303=>x"00133",
4304=>x"00133",
4305=>x"00133",
4306=>x"00133",
4307=>x"00133",
4308=>x"00133",
4309=>x"00133",
4310=>x"00133",
4311=>x"00133",
4312=>x"00134",
4313=>x"00134",
4314=>x"00134",
4315=>x"00134",
4316=>x"00134",
4317=>x"00134",
4318=>x"00134",
4319=>x"00134",
4320=>x"00134",
4321=>x"00134",
4322=>x"00134",
4323=>x"00134",
4324=>x"00134",
4325=>x"00134",
4326=>x"00135",
4327=>x"00135",
4328=>x"00135",
4329=>x"00135",
4330=>x"00135",
4331=>x"00135",
4332=>x"00135",
4333=>x"00135",
4334=>x"00135",
4335=>x"00135",
4336=>x"00135",
4337=>x"00135",
4338=>x"00135",
4339=>x"00135",
4340=>x"00136",
4341=>x"00136",
4342=>x"00136",
4343=>x"00136",
4344=>x"00136",
4345=>x"00136",
4346=>x"00136",
4347=>x"00136",
4348=>x"00136",
4349=>x"00136",
4350=>x"00136",
4351=>x"00136",
4352=>x"00136",
4353=>x"00136",
4354=>x"00137",
4355=>x"00137",
4356=>x"00137",
4357=>x"00137",
4358=>x"00137",
4359=>x"00137",
4360=>x"00137",
4361=>x"00137",
4362=>x"00137",
4363=>x"00137",
4364=>x"00137",
4365=>x"00137",
4366=>x"00137",
4367=>x"00137",
4368=>x"00138",
4369=>x"00138",
4370=>x"00138",
4371=>x"00138",
4372=>x"00138",
4373=>x"00138",
4374=>x"00138",
4375=>x"00138",
4376=>x"00138",
4377=>x"00138",
4378=>x"00138",
4379=>x"00138",
4380=>x"00138",
4381=>x"00138",
4382=>x"00139",
4383=>x"00139",
4384=>x"00139",
4385=>x"00139",
4386=>x"00139",
4387=>x"00139",
4388=>x"00139",
4389=>x"00139",
4390=>x"00139",
4391=>x"00139",
4392=>x"00139",
4393=>x"00139",
4394=>x"00139",
4395=>x"00139",
4396=>x"0013a",
4397=>x"0013a",
4398=>x"0013a",
4399=>x"0013a",
4400=>x"0013a",
4401=>x"0013a",
4402=>x"0013a",
4403=>x"0013a",
4404=>x"0013a",
4405=>x"0013a",
4406=>x"0013a",
4407=>x"0013a",
4408=>x"0013a",
4409=>x"0013a",
4410=>x"0013b",
4411=>x"0013b",
4412=>x"0013b",
4413=>x"0013b",
4414=>x"0013b",
4415=>x"0013b",
4416=>x"0013b",
4417=>x"0013b",
4418=>x"0013b",
4419=>x"0013b",
4420=>x"0013b",
4421=>x"0013b",
4422=>x"0013b",
4423=>x"0013b",
4424=>x"0013c",
4425=>x"0013c",
4426=>x"0013c",
4427=>x"0013c",
4428=>x"0013c",
4429=>x"0013c",
4430=>x"0013c",
4431=>x"0013c",
4432=>x"0013c",
4433=>x"0013c",
4434=>x"0013c",
4435=>x"0013c",
4436=>x"0013c",
4437=>x"0013c",
4438=>x"0013d",
4439=>x"0013d",
4440=>x"0013d",
4441=>x"0013d",
4442=>x"0013d",
4443=>x"0013d",
4444=>x"0013d",
4445=>x"0013d",
4446=>x"0013d",
4447=>x"0013d",
4448=>x"0013d",
4449=>x"0013d",
4450=>x"0013d",
4451=>x"0013d",
4452=>x"0013e",
4453=>x"0013e",
4454=>x"0013e",
4455=>x"0013e",
4456=>x"0013e",
4457=>x"0013e",
4458=>x"0013e",
4459=>x"0013e",
4460=>x"0013e",
4461=>x"0013e",
4462=>x"0013e",
4463=>x"0013e",
4464=>x"0013e",
4465=>x"0013e",
4466=>x"0013f",
4467=>x"0013f",
4468=>x"0013f",
4469=>x"0013f",
4470=>x"0013f",
4471=>x"0013f",
4472=>x"0013f",
4473=>x"0013f",
4474=>x"0013f",
4475=>x"0013f",
4476=>x"0013f",
4477=>x"0013f",
4478=>x"0013f",
4479=>x"0013f",
4480=>x"00140",
4481=>x"00140",
4482=>x"00140",
4483=>x"00140",
4484=>x"00140",
4485=>x"00140",
4486=>x"00140",
4487=>x"00140",
4488=>x"00140",
4489=>x"00140",
4490=>x"00140",
4491=>x"00140",
4492=>x"00140",
4493=>x"00140",
4494=>x"00141",
4495=>x"00141",
4496=>x"00141",
4497=>x"00141",
4498=>x"00141",
4499=>x"00141",
4500=>x"00141",
4501=>x"00141",
4502=>x"00141",
4503=>x"00141",
4504=>x"00141",
4505=>x"00141",
4506=>x"00141",
4507=>x"00141",
4508=>x"00142",
4509=>x"00142",
4510=>x"00142",
4511=>x"00142",
4512=>x"00142",
4513=>x"00142",
4514=>x"00142",
4515=>x"00142",
4516=>x"00142",
4517=>x"00142",
4518=>x"00142",
4519=>x"00142",
4520=>x"00142",
4521=>x"00142",
4522=>x"00143",
4523=>x"00143",
4524=>x"00143",
4525=>x"00143",
4526=>x"00143",
4527=>x"00143",
4528=>x"00143",
4529=>x"00143",
4530=>x"00143",
4531=>x"00143",
4532=>x"00143",
4533=>x"00143",
4534=>x"00143",
4535=>x"00143",
4536=>x"00144",
4537=>x"00144",
4538=>x"00144",
4539=>x"00144",
4540=>x"00144",
4541=>x"00144",
4542=>x"00144",
4543=>x"00144",
4544=>x"00144",
4545=>x"00144",
4546=>x"00144",
4547=>x"00144",
4548=>x"00144",
4549=>x"00144",
4550=>x"00145",
4551=>x"00145",
4552=>x"00145",
4553=>x"00145",
4554=>x"00145",
4555=>x"00145",
4556=>x"00145",
4557=>x"00145",
4558=>x"00145",
4559=>x"00145",
4560=>x"00145",
4561=>x"00145",
4562=>x"00145",
4563=>x"00145",
4564=>x"00146",
4565=>x"00146",
4566=>x"00146",
4567=>x"00146",
4568=>x"00146",
4569=>x"00146",
4570=>x"00146",
4571=>x"00146",
4572=>x"00146",
4573=>x"00146",
4574=>x"00146",
4575=>x"00146",
4576=>x"00146",
4577=>x"00146",
4578=>x"00147",
4579=>x"00147",
4580=>x"00147",
4581=>x"00147",
4582=>x"00147",
4583=>x"00147",
4584=>x"00147",
4585=>x"00147",
4586=>x"00147",
4587=>x"00147",
4588=>x"00147",
4589=>x"00147",
4590=>x"00147",
4591=>x"00147",
4592=>x"00148",
4593=>x"00148",
4594=>x"00148",
4595=>x"00148",
4596=>x"00148",
4597=>x"00148",
4598=>x"00148",
4599=>x"00148",
4600=>x"00148",
4601=>x"00148",
4602=>x"00148",
4603=>x"00148",
4604=>x"00148",
4605=>x"00148",
4606=>x"00149",
4607=>x"00149",
4608=>x"00149",
4609=>x"00149",
4610=>x"00149",
4611=>x"00149",
4612=>x"00149",
4613=>x"00149",
4614=>x"00149",
4615=>x"00149",
4616=>x"00149",
4617=>x"00149",
4618=>x"00149",
4619=>x"00149",
4620=>x"0014a",
4621=>x"0014a",
4622=>x"0014a",
4623=>x"0014a",
4624=>x"0014a",
4625=>x"0014a",
4626=>x"0014a",
4627=>x"0014a",
4628=>x"0014a",
4629=>x"0014a",
4630=>x"0014a",
4631=>x"0014a",
4632=>x"0014a",
4633=>x"0014a",
4634=>x"0014b",
4635=>x"0014b",
4636=>x"0014b",
4637=>x"0014b",
4638=>x"0014b",
4639=>x"0014b",
4640=>x"0014b",
4641=>x"0014b",
4642=>x"0014b",
4643=>x"0014b",
4644=>x"0014b",
4645=>x"0014b",
4646=>x"0014b",
4647=>x"0014b",
4648=>x"0014c",
4649=>x"0014c",
4650=>x"0014c",
4651=>x"0014c",
4652=>x"0014c",
4653=>x"0014c",
4654=>x"0014c",
4655=>x"0014c",
4656=>x"0014c",
4657=>x"0014c",
4658=>x"0014c",
4659=>x"0014c",
4660=>x"0014c",
4661=>x"0014c",
4662=>x"0014d",
4663=>x"0014d",
4664=>x"0014d",
4665=>x"0014d",
4666=>x"0014d",
4667=>x"0014d",
4668=>x"0014d",
4669=>x"0014d",
4670=>x"0014d",
4671=>x"0014d",
4672=>x"0014d",
4673=>x"0014d",
4674=>x"0014d",
4675=>x"0014d",
4676=>x"0014e",
4677=>x"0014e",
4678=>x"0014e",
4679=>x"0014e",
4680=>x"0014e",
4681=>x"0014e",
4682=>x"0014e",
4683=>x"0014e",
4684=>x"0014e",
4685=>x"0014e",
4686=>x"0014e",
4687=>x"0014e",
4688=>x"0014e",
4689=>x"0014e",
4690=>x"0014f",
4691=>x"0014f",
4692=>x"0014f",
4693=>x"0014f",
4694=>x"0014f",
4695=>x"0014f",
4696=>x"0014f",
4697=>x"0014f",
4698=>x"0014f",
4699=>x"0014f",
4700=>x"0014f",
4701=>x"0014f",
4702=>x"0014f",
4703=>x"0014f",
4704=>x"00150",
4705=>x"00150",
4706=>x"00150",
4707=>x"00150",
4708=>x"00150",
4709=>x"00150",
4710=>x"00150",
4711=>x"00150",
4712=>x"00150",
4713=>x"00150",
4714=>x"00150",
4715=>x"00150",
4716=>x"00150",
4717=>x"00150",
4718=>x"00151",
4719=>x"00151",
4720=>x"00151",
4721=>x"00151",
4722=>x"00151",
4723=>x"00151",
4724=>x"00151",
4725=>x"00151",
4726=>x"00151",
4727=>x"00151",
4728=>x"00151",
4729=>x"00151",
4730=>x"00151",
4731=>x"00151",
4732=>x"00152",
4733=>x"00152",
4734=>x"00152",
4735=>x"00152",
4736=>x"00152",
4737=>x"00152",
4738=>x"00152",
4739=>x"00152",
4740=>x"00152",
4741=>x"00152",
4742=>x"00152",
4743=>x"00152",
4744=>x"00152",
4745=>x"00152",
4746=>x"00153",
4747=>x"00153",
4748=>x"00153",
4749=>x"00153",
4750=>x"00153",
4751=>x"00153",
4752=>x"00153",
4753=>x"00153",
4754=>x"00153",
4755=>x"00153",
4756=>x"00153",
4757=>x"00153",
4758=>x"00153",
4759=>x"00153",
4760=>x"00154",
4761=>x"00154",
4762=>x"00154",
4763=>x"00154",
4764=>x"00154",
4765=>x"00154",
4766=>x"00154",
4767=>x"00154",
4768=>x"00154",
4769=>x"00154",
4770=>x"00154",
4771=>x"00154",
4772=>x"00154",
4773=>x"00154",
4774=>x"00155",
4775=>x"00155",
4776=>x"00155",
4777=>x"00155",
4778=>x"00155",
4779=>x"00155",
4780=>x"00155",
4781=>x"00155",
4782=>x"00155",
4783=>x"00155",
4784=>x"00155",
4785=>x"00155",
4786=>x"00155",
4787=>x"00155",
4788=>x"00156",
4789=>x"00156",
4790=>x"00156",
4791=>x"00156",
4792=>x"00156",
4793=>x"00156",
4794=>x"00156",
4795=>x"00156",
4796=>x"00156",
4797=>x"00156",
4798=>x"00156",
4799=>x"00156",
4800=>x"00156",
4801=>x"00156",
4802=>x"00157",
4803=>x"00157",
4804=>x"00157",
4805=>x"00157",
4806=>x"00157",
4807=>x"00157",
4808=>x"00157",
4809=>x"00157",
4810=>x"00157",
4811=>x"00157",
4812=>x"00157",
4813=>x"00157",
4814=>x"00157",
4815=>x"00157",
4816=>x"00158",
4817=>x"00158",
4818=>x"00158",
4819=>x"00158",
4820=>x"00158",
4821=>x"00158",
4822=>x"00158",
4823=>x"00158",
4824=>x"00158",
4825=>x"00158",
4826=>x"00158",
4827=>x"00158",
4828=>x"00158",
4829=>x"00158",
4830=>x"00159",
4831=>x"00159",
4832=>x"00159",
4833=>x"00159",
4834=>x"00159",
4835=>x"00159",
4836=>x"00159",
4837=>x"00159",
4838=>x"00159",
4839=>x"00159",
4840=>x"00159",
4841=>x"00159",
4842=>x"00159",
4843=>x"00159",
4844=>x"0015a",
4845=>x"0015a",
4846=>x"0015a",
4847=>x"0015a",
4848=>x"0015a",
4849=>x"0015a",
4850=>x"0015a",
4851=>x"0015a",
4852=>x"0015a",
4853=>x"0015a",
4854=>x"0015a",
4855=>x"0015a",
4856=>x"0015a",
4857=>x"0015a",
4858=>x"0015b",
4859=>x"0015b",
4860=>x"0015b",
4861=>x"0015b",
4862=>x"0015b",
4863=>x"0015b",
4864=>x"0015b",
4865=>x"0015b",
4866=>x"0015b",
4867=>x"0015b",
4868=>x"0015b",
4869=>x"0015b",
4870=>x"0015b",
4871=>x"0015b",
4872=>x"0015c",
4873=>x"0015c",
4874=>x"0015c",
4875=>x"0015c",
4876=>x"0015c",
4877=>x"0015c",
4878=>x"0015c",
4879=>x"0015c",
4880=>x"0015c",
4881=>x"0015c",
4882=>x"0015c",
4883=>x"0015c",
4884=>x"0015c",
4885=>x"0015c",
4886=>x"0015d",
4887=>x"0015d",
4888=>x"0015d",
4889=>x"0015d",
4890=>x"0015d",
4891=>x"0015d",
4892=>x"0015d",
4893=>x"0015d",
4894=>x"0015d",
4895=>x"0015d",
4896=>x"0015d",
4897=>x"0015d",
4898=>x"0015d",
4899=>x"0015d",
4900=>x"0015e",
4901=>x"0015e",
4902=>x"0015e",
4903=>x"0015e",
4904=>x"0015e",
4905=>x"0015e",
4906=>x"0015e",
4907=>x"0015e",
4908=>x"0015e",
4909=>x"0015e",
4910=>x"0015e",
4911=>x"0015e",
4912=>x"0015e",
4913=>x"0015e",
4914=>x"0015f",
4915=>x"0015f",
4916=>x"0015f",
4917=>x"0015f",
4918=>x"0015f",
4919=>x"0015f",
4920=>x"0015f",
4921=>x"0015f",
4922=>x"0015f",
4923=>x"0015f",
4924=>x"0015f",
4925=>x"0015f",
4926=>x"0015f",
4927=>x"0015f",
4928=>x"00160",
4929=>x"00160",
4930=>x"00160",
4931=>x"00160",
4932=>x"00160",
4933=>x"00160",
4934=>x"00160",
4935=>x"00160",
4936=>x"00160",
4937=>x"00160",
4938=>x"00160",
4939=>x"00160",
4940=>x"00160",
4941=>x"00160",
4942=>x"00161",
4943=>x"00161",
4944=>x"00161",
4945=>x"00161",
4946=>x"00161",
4947=>x"00161",
4948=>x"00161",
4949=>x"00161",
4950=>x"00161",
4951=>x"00161",
4952=>x"00161",
4953=>x"00161",
4954=>x"00161",
4955=>x"00161",
4956=>x"00162",
4957=>x"00162",
4958=>x"00162",
4959=>x"00162",
4960=>x"00162",
4961=>x"00162",
4962=>x"00162",
4963=>x"00162",
4964=>x"00162",
4965=>x"00162",
4966=>x"00162",
4967=>x"00162",
4968=>x"00162",
4969=>x"00162",
4970=>x"00163",
4971=>x"00163",
4972=>x"00163",
4973=>x"00163",
4974=>x"00163",
4975=>x"00163",
4976=>x"00163",
4977=>x"00163",
4978=>x"00163",
4979=>x"00163",
4980=>x"00163",
4981=>x"00163",
4982=>x"00163",
4983=>x"00163",
4984=>x"00164",
4985=>x"00164",
4986=>x"00164",
4987=>x"00164",
4988=>x"00164",
4989=>x"00164",
4990=>x"00164",
4991=>x"00164",
4992=>x"00164",
4993=>x"00164",
4994=>x"00164",
4995=>x"00164",
4996=>x"00164",
4997=>x"00164",
4998=>x"00165",
4999=>x"00165",
5000=>x"00165",
5001=>x"00165",
5002=>x"00165",
5003=>x"00165",
5004=>x"00165",
5005=>x"00165",
5006=>x"00165",
5007=>x"00165",
5008=>x"00165",
5009=>x"00165",
5010=>x"00165",
5011=>x"00165",
5012=>x"00166",
5013=>x"00166",
5014=>x"00166",
5015=>x"00166",
5016=>x"00166",
5017=>x"00166",
5018=>x"00166",
5019=>x"00166",
5020=>x"00166",
5021=>x"00166",
5022=>x"00166",
5023=>x"00166",
5024=>x"00166",
5025=>x"00166",
5026=>x"00167",
5027=>x"00167",
5028=>x"00167",
5029=>x"00167",
5030=>x"00167",
5031=>x"00167",
5032=>x"00167",
5033=>x"00167",
5034=>x"00167",
5035=>x"00167",
5036=>x"00167",
5037=>x"00167",
5038=>x"00167",
5039=>x"00167",
5040=>x"00168",
5041=>x"00168",
5042=>x"00168",
5043=>x"00168",
5044=>x"00168",
5045=>x"00168",
5046=>x"00168",
5047=>x"00168",
5048=>x"00168",
5049=>x"00168",
5050=>x"00168",
5051=>x"00168",
5052=>x"00168",
5053=>x"00168",
5054=>x"00169",
5055=>x"00169",
5056=>x"00169",
5057=>x"00169",
5058=>x"00169",
5059=>x"00169",
5060=>x"00169",
5061=>x"00169",
5062=>x"00169",
5063=>x"00169",
5064=>x"00169",
5065=>x"00169",
5066=>x"00169",
5067=>x"00169",
5068=>x"0016a",
5069=>x"0016a",
5070=>x"0016a",
5071=>x"0016a",
5072=>x"0016a",
5073=>x"0016a",
5074=>x"0016a",
5075=>x"0016a",
5076=>x"0016a",
5077=>x"0016a",
5078=>x"0016a",
5079=>x"0016a",
5080=>x"0016a",
5081=>x"0016a",
5082=>x"0016b",
5083=>x"0016b",
5084=>x"0016b",
5085=>x"0016b",
5086=>x"0016b",
5087=>x"0016b",
5088=>x"0016b",
5089=>x"0016b",
5090=>x"0016b",
5091=>x"0016b",
5092=>x"0016b",
5093=>x"0016b",
5094=>x"0016b",
5095=>x"0016b",
5096=>x"0016c",
5097=>x"0016c",
5098=>x"0016c",
5099=>x"0016c",
5100=>x"0016c",
5101=>x"0016c",
5102=>x"0016c",
5103=>x"0016c",
5104=>x"0016c",
5105=>x"0016c",
5106=>x"0016c",
5107=>x"0016c",
5108=>x"0016c",
5109=>x"0016c",
5110=>x"0016d",
5111=>x"0016d",
5112=>x"0016d",
5113=>x"0016d",
5114=>x"0016d",
5115=>x"0016d",
5116=>x"0016d",
5117=>x"0016d",
5118=>x"0016d",
5119=>x"0016d",
5120=>x"0016d",
5121=>x"0016d",
5122=>x"0016d",
5123=>x"0016d",
5124=>x"0016e",
5125=>x"0016e",
5126=>x"0016e",
5127=>x"0016e",
5128=>x"0016e",
5129=>x"0016e",
5130=>x"0016e",
5131=>x"0016e",
5132=>x"0016e",
5133=>x"0016e",
5134=>x"0016e",
5135=>x"0016e",
5136=>x"0016e",
5137=>x"0016e",
5138=>x"0016f",
5139=>x"0016f",
5140=>x"0016f",
5141=>x"0016f",
5142=>x"0016f",
5143=>x"0016f",
5144=>x"0016f",
5145=>x"0016f",
5146=>x"0016f",
5147=>x"0016f",
5148=>x"0016f",
5149=>x"0016f",
5150=>x"0016f",
5151=>x"0016f",
5152=>x"00170",
5153=>x"00170",
5154=>x"00170",
5155=>x"00170",
5156=>x"00170",
5157=>x"00170",
5158=>x"00170",
5159=>x"00170",
5160=>x"00170",
5161=>x"00170",
5162=>x"00170",
5163=>x"00170",
5164=>x"00170",
5165=>x"00170",
5166=>x"00171",
5167=>x"00171",
5168=>x"00171",
5169=>x"00171",
5170=>x"00171",
5171=>x"00171",
5172=>x"00171",
5173=>x"00171",
5174=>x"00171",
5175=>x"00171",
5176=>x"00171",
5177=>x"00171",
5178=>x"00171",
5179=>x"00171",
5180=>x"00172",
5181=>x"00172",
5182=>x"00172",
5183=>x"00172",
5184=>x"00172",
5185=>x"00172",
5186=>x"00172",
5187=>x"00172",
5188=>x"00172",
5189=>x"00172",
5190=>x"00172",
5191=>x"00172",
5192=>x"00172",
5193=>x"00172",
5194=>x"00173",
5195=>x"00173",
5196=>x"00173",
5197=>x"00173",
5198=>x"00173",
5199=>x"00173",
5200=>x"00173",
5201=>x"00173",
5202=>x"00173",
5203=>x"00173",
5204=>x"00173",
5205=>x"00173",
5206=>x"00173",
5207=>x"00173",
5208=>x"00174",
5209=>x"00174",
5210=>x"00174",
5211=>x"00174",
5212=>x"00174",
5213=>x"00174",
5214=>x"00174",
5215=>x"00174",
5216=>x"00174",
5217=>x"00174",
5218=>x"00174",
5219=>x"00174",
5220=>x"00174",
5221=>x"00174",
5222=>x"00175",
5223=>x"00175",
5224=>x"00175",
5225=>x"00175",
5226=>x"00175",
5227=>x"00175",
5228=>x"00175",
5229=>x"00175",
5230=>x"00175",
5231=>x"00175",
5232=>x"00175",
5233=>x"00175",
5234=>x"00175",
5235=>x"00175",
5236=>x"00176",
5237=>x"00176",
5238=>x"00176",
5239=>x"00176",
5240=>x"00176",
5241=>x"00176",
5242=>x"00176",
5243=>x"00176",
5244=>x"00176",
5245=>x"00176",
5246=>x"00176",
5247=>x"00176",
5248=>x"00176",
5249=>x"00176",
5250=>x"00177",
5251=>x"00177",
5252=>x"00177",
5253=>x"00177",
5254=>x"00177",
5255=>x"00177",
5256=>x"00177",
5257=>x"00177",
5258=>x"00177",
5259=>x"00177",
5260=>x"00177",
5261=>x"00177",
5262=>x"00177",
5263=>x"00177",
5264=>x"00178",
5265=>x"00178",
5266=>x"00178",
5267=>x"00178",
5268=>x"00178",
5269=>x"00178",
5270=>x"00178",
5271=>x"00178",
5272=>x"00178",
5273=>x"00178",
5274=>x"00178",
5275=>x"00178",
5276=>x"00178",
5277=>x"00178",
5278=>x"00179",
5279=>x"00179",
5280=>x"00179",
5281=>x"00179",
5282=>x"00179",
5283=>x"00179",
5284=>x"00179",
5285=>x"00179",
5286=>x"00179",
5287=>x"00179",
5288=>x"00179",
5289=>x"00179",
5290=>x"00179",
5291=>x"00179",
5292=>x"0017a",
5293=>x"0017a",
5294=>x"0017a",
5295=>x"0017a",
5296=>x"0017a",
5297=>x"0017a",
5298=>x"0017a",
5299=>x"0017a",
5300=>x"0017a",
5301=>x"0017a",
5302=>x"0017a",
5303=>x"0017a",
5304=>x"0017a",
5305=>x"0017a",
5306=>x"0017b",
5307=>x"0017b",
5308=>x"0017b",
5309=>x"0017b",
5310=>x"0017b",
5311=>x"0017b",
5312=>x"0017b",
5313=>x"0017b",
5314=>x"0017b",
5315=>x"0017b",
5316=>x"0017b",
5317=>x"0017b",
5318=>x"0017b",
5319=>x"0017b",
5320=>x"0017c",
5321=>x"0017c",
5322=>x"0017c",
5323=>x"0017c",
5324=>x"0017c",
5325=>x"0017c",
5326=>x"0017c",
5327=>x"0017c",
5328=>x"0017c",
5329=>x"0017c",
5330=>x"0017c",
5331=>x"0017c",
5332=>x"0017c",
5333=>x"0017c",
5334=>x"0017d",
5335=>x"0017d",
5336=>x"0017d",
5337=>x"0017d",
5338=>x"0017d",
5339=>x"0017d",
5340=>x"0017d",
5341=>x"0017d",
5342=>x"0017d",
5343=>x"0017d",
5344=>x"0017d",
5345=>x"0017d",
5346=>x"0017d",
5347=>x"0017d",
5348=>x"0017e",
5349=>x"0017e",
5350=>x"0017e",
5351=>x"0017e",
5352=>x"0017e",
5353=>x"0017e",
5354=>x"0017e",
5355=>x"0017e",
5356=>x"0017e",
5357=>x"0017e",
5358=>x"0017e",
5359=>x"0017e",
5360=>x"0017e",
5361=>x"0017e",
5362=>x"0017f",
5363=>x"0017f",
5364=>x"0017f",
5365=>x"0017f",
5366=>x"0017f",
5367=>x"0017f",
5368=>x"0017f",
5369=>x"0017f",
5370=>x"0017f",
5371=>x"0017f",
5372=>x"0017f",
5373=>x"0017f",
5374=>x"0017f",
5375=>x"0017f",
5376=>x"00180",
5377=>x"00180",
5378=>x"00180",
5379=>x"00180",
5380=>x"00180",
5381=>x"00180",
5382=>x"00180",
5383=>x"00180",
5384=>x"00180",
5385=>x"00180",
5386=>x"00180",
5387=>x"00180",
5388=>x"00180",
5389=>x"00180",
5390=>x"00181",
5391=>x"00181",
5392=>x"00181",
5393=>x"00181",
5394=>x"00181",
5395=>x"00181",
5396=>x"00181",
5397=>x"00181",
5398=>x"00181",
5399=>x"00181",
5400=>x"00181",
5401=>x"00181",
5402=>x"00181",
5403=>x"00181",
5404=>x"00182",
5405=>x"00182",
5406=>x"00182",
5407=>x"00182",
5408=>x"00182",
5409=>x"00182",
5410=>x"00182",
5411=>x"00182",
5412=>x"00182",
5413=>x"00182",
5414=>x"00182",
5415=>x"00182",
5416=>x"00182",
5417=>x"00182",
5418=>x"00183",
5419=>x"00183",
5420=>x"00183",
5421=>x"00183",
5422=>x"00183",
5423=>x"00183",
5424=>x"00183",
5425=>x"00183",
5426=>x"00183",
5427=>x"00183",
5428=>x"00183",
5429=>x"00183",
5430=>x"00183",
5431=>x"00183",
5432=>x"00184",
5433=>x"00184",
5434=>x"00184",
5435=>x"00184",
5436=>x"00184",
5437=>x"00184",
5438=>x"00184",
5439=>x"00184",
5440=>x"00184",
5441=>x"00184",
5442=>x"00184",
5443=>x"00184",
5444=>x"00184",
5445=>x"00184",
5446=>x"00185",
5447=>x"00185",
5448=>x"00185",
5449=>x"00185",
5450=>x"00185",
5451=>x"00185",
5452=>x"00185",
5453=>x"00185",
5454=>x"00185",
5455=>x"00185",
5456=>x"00185",
5457=>x"00185",
5458=>x"00185",
5459=>x"00185",
5460=>x"00186",
5461=>x"00186",
5462=>x"00186",
5463=>x"00186",
5464=>x"00186",
5465=>x"00186",
5466=>x"00186",
5467=>x"00186",
5468=>x"00186",
5469=>x"00186",
5470=>x"00186",
5471=>x"00186",
5472=>x"00186",
5473=>x"00186",
5474=>x"00187",
5475=>x"00187",
5476=>x"00187",
5477=>x"00187",
5478=>x"00187",
5479=>x"00187",
5480=>x"00187",
5481=>x"00187",
5482=>x"00187",
5483=>x"00187",
5484=>x"00187",
5485=>x"00187",
5486=>x"00187",
5487=>x"00187",
5488=>x"00188",
5489=>x"00188",
5490=>x"00188",
5491=>x"00188",
5492=>x"00188",
5493=>x"00188",
5494=>x"00188",
5495=>x"00188",
5496=>x"00188",
5497=>x"00188",
5498=>x"00188",
5499=>x"00188",
5500=>x"00188",
5501=>x"00188",
5502=>x"00189",
5503=>x"00189",
5504=>x"00189",
5505=>x"00189",
5506=>x"00189",
5507=>x"00189",
5508=>x"00189",
5509=>x"00189",
5510=>x"00189",
5511=>x"00189",
5512=>x"00189",
5513=>x"00189",
5514=>x"00189",
5515=>x"00189",
5516=>x"0018a",
5517=>x"0018a",
5518=>x"0018a",
5519=>x"0018a",
5520=>x"0018a",
5521=>x"0018a",
5522=>x"0018a",
5523=>x"0018a",
5524=>x"0018a",
5525=>x"0018a",
5526=>x"0018a",
5527=>x"0018a",
5528=>x"0018a",
5529=>x"0018a",
5530=>x"0018b",
5531=>x"0018b",
5532=>x"0018b",
5533=>x"0018b",
5534=>x"0018b",
5535=>x"0018b",
5536=>x"0018b",
5537=>x"0018b",
5538=>x"0018b",
5539=>x"0018b",
5540=>x"0018b",
5541=>x"0018b",
5542=>x"0018b",
5543=>x"0018b",
5544=>x"0018c",
5545=>x"0018c",
5546=>x"0018c",
5547=>x"0018c",
5548=>x"0018c",
5549=>x"0018c",
5550=>x"0018c",
5551=>x"0018c",
5552=>x"0018c",
5553=>x"0018c",
5554=>x"0018c",
5555=>x"0018c",
5556=>x"0018c",
5557=>x"0018c",
5558=>x"0018d",
5559=>x"0018d",
5560=>x"0018d",
5561=>x"0018d",
5562=>x"0018d",
5563=>x"0018d",
5564=>x"0018d",
5565=>x"0018d",
5566=>x"0018d",
5567=>x"0018d",
5568=>x"0018d",
5569=>x"0018d",
5570=>x"0018d",
5571=>x"0018d",
5572=>x"0018e",
5573=>x"0018e",
5574=>x"0018e",
5575=>x"0018e",
5576=>x"0018e",
5577=>x"0018e",
5578=>x"0018e",
5579=>x"0018e",
5580=>x"0018e",
5581=>x"0018e",
5582=>x"0018e",
5583=>x"0018e",
5584=>x"0018e",
5585=>x"0018e",
5586=>x"0018f",
5587=>x"0018f",
5588=>x"0018f",
5589=>x"0018f",
5590=>x"0018f",
5591=>x"0018f",
5592=>x"0018f",
5593=>x"0018f",
5594=>x"0018f",
5595=>x"0018f",
5596=>x"0018f",
5597=>x"0018f",
5598=>x"0018f",
5599=>x"0018f",
5600=>x"00190",
5601=>x"00190",
5602=>x"00190",
5603=>x"00190",
5604=>x"00190",
5605=>x"00190",
5606=>x"00190",
5607=>x"00190",
5608=>x"00190",
5609=>x"00190",
5610=>x"00190",
5611=>x"00190",
5612=>x"00190",
5613=>x"00190",
5614=>x"00191",
5615=>x"00191",
5616=>x"00191",
5617=>x"00191",
5618=>x"00191",
5619=>x"00191",
5620=>x"00191",
5621=>x"00191",
5622=>x"00191",
5623=>x"00191",
5624=>x"00191",
5625=>x"00191",
5626=>x"00191",
5627=>x"00191",
5628=>x"00192",
5629=>x"00192",
5630=>x"00192",
5631=>x"00192",
5632=>x"00192",
5633=>x"00192",
5634=>x"00192",
5635=>x"00192",
5636=>x"00192",
5637=>x"00192",
5638=>x"00192",
5639=>x"00192",
5640=>x"00192",
5641=>x"00192",
5642=>x"00193",
5643=>x"00193",
5644=>x"00193",
5645=>x"00193",
5646=>x"00193",
5647=>x"00193",
5648=>x"00193",
5649=>x"00193",
5650=>x"00193",
5651=>x"00193",
5652=>x"00193",
5653=>x"00193",
5654=>x"00193",
5655=>x"00193",
5656=>x"00194",
5657=>x"00194",
5658=>x"00194",
5659=>x"00194",
5660=>x"00194",
5661=>x"00194",
5662=>x"00194",
5663=>x"00194",
5664=>x"00194",
5665=>x"00194",
5666=>x"00194",
5667=>x"00194",
5668=>x"00194",
5669=>x"00194",
5670=>x"00195",
5671=>x"00195",
5672=>x"00195",
5673=>x"00195",
5674=>x"00195",
5675=>x"00195",
5676=>x"00195",
5677=>x"00195",
5678=>x"00195",
5679=>x"00195",
5680=>x"00195",
5681=>x"00195",
5682=>x"00195",
5683=>x"00195",
5684=>x"00196",
5685=>x"00196",
5686=>x"00196",
5687=>x"00196",
5688=>x"00196",
5689=>x"00196",
5690=>x"00196",
5691=>x"00196",
5692=>x"00196",
5693=>x"00196",
5694=>x"00196",
5695=>x"00196",
5696=>x"00196",
5697=>x"00196",
5698=>x"00197",
5699=>x"00197",
5700=>x"00197",
5701=>x"00197",
5702=>x"00197",
5703=>x"00197",
5704=>x"00197",
5705=>x"00197",
5706=>x"00197",
5707=>x"00197",
5708=>x"00197",
5709=>x"00197",
5710=>x"00197",
5711=>x"00197",
5712=>x"00198",
5713=>x"00198",
5714=>x"00198",
5715=>x"00198",
5716=>x"00198",
5717=>x"00198",
5718=>x"00198",
5719=>x"00198",
5720=>x"00198",
5721=>x"00198",
5722=>x"00198",
5723=>x"00198",
5724=>x"00198",
5725=>x"00198",
5726=>x"00199",
5727=>x"00199",
5728=>x"00199",
5729=>x"00199",
5730=>x"00199",
5731=>x"00199",
5732=>x"00199",
5733=>x"00199",
5734=>x"00199",
5735=>x"00199",
5736=>x"00199",
5737=>x"00199",
5738=>x"00199",
5739=>x"00199",
5740=>x"0019a",
5741=>x"0019a",
5742=>x"0019a",
5743=>x"0019a",
5744=>x"0019a",
5745=>x"0019a",
5746=>x"0019a",
5747=>x"0019a",
5748=>x"0019a",
5749=>x"0019a",
5750=>x"0019a",
5751=>x"0019a",
5752=>x"0019a",
5753=>x"0019a",
5754=>x"0019b",
5755=>x"0019b",
5756=>x"0019b",
5757=>x"0019b",
5758=>x"0019b",
5759=>x"0019b",
5760=>x"0019b",
5761=>x"0019b",
5762=>x"0019b",
5763=>x"0019b",
5764=>x"0019b",
5765=>x"0019b",
5766=>x"0019b",
5767=>x"0019b",
5768=>x"0019c",
5769=>x"0019c",
5770=>x"0019c",
5771=>x"0019c",
5772=>x"0019c",
5773=>x"0019c",
5774=>x"0019c",
5775=>x"0019c",
5776=>x"0019c",
5777=>x"0019c",
5778=>x"0019c",
5779=>x"0019c",
5780=>x"0019c",
5781=>x"0019c",
5782=>x"0019d",
5783=>x"0019d",
5784=>x"0019d",
5785=>x"0019d",
5786=>x"0019d",
5787=>x"0019d",
5788=>x"0019d",
5789=>x"0019d",
5790=>x"0019d",
5791=>x"0019d",
5792=>x"0019d",
5793=>x"0019d",
5794=>x"0019d",
5795=>x"0019d",
5796=>x"0019e",
5797=>x"0019e",
5798=>x"0019e",
5799=>x"0019e",
5800=>x"0019e",
5801=>x"0019e",
5802=>x"0019e",
5803=>x"0019e",
5804=>x"0019e",
5805=>x"0019e",
5806=>x"0019e",
5807=>x"0019e",
5808=>x"0019e",
5809=>x"0019e",
5810=>x"0019f",
5811=>x"0019f",
5812=>x"0019f",
5813=>x"0019f",
5814=>x"0019f",
5815=>x"0019f",
5816=>x"0019f",
5817=>x"0019f",
5818=>x"0019f",
5819=>x"0019f",
5820=>x"0019f",
5821=>x"0019f",
5822=>x"0019f",
5823=>x"0019f",
5824=>x"001a0",
5825=>x"001a0",
5826=>x"001a0",
5827=>x"001a0",
5828=>x"001a0",
5829=>x"001a0",
5830=>x"001a0",
5831=>x"001a0",
5832=>x"001a0",
5833=>x"001a0",
5834=>x"001a0",
5835=>x"001a0",
5836=>x"001a0",
5837=>x"001a0",
5838=>x"001a1",
5839=>x"001a1",
5840=>x"001a1",
5841=>x"001a1",
5842=>x"001a1",
5843=>x"001a1",
5844=>x"001a1",
5845=>x"001a1",
5846=>x"001a1",
5847=>x"001a1",
5848=>x"001a1",
5849=>x"001a1",
5850=>x"001a1",
5851=>x"001a1",
5852=>x"001a2",
5853=>x"001a2",
5854=>x"001a2",
5855=>x"001a2",
5856=>x"001a2",
5857=>x"001a2",
5858=>x"001a2",
5859=>x"001a2",
5860=>x"001a2",
5861=>x"001a2",
5862=>x"001a2",
5863=>x"001a2",
5864=>x"001a2",
5865=>x"001a2",
5866=>x"001a3",
5867=>x"001a3",
5868=>x"001a3",
5869=>x"001a3",
5870=>x"001a3",
5871=>x"001a3",
5872=>x"001a3",
5873=>x"001a3",
5874=>x"001a3",
5875=>x"001a3",
5876=>x"001a3",
5877=>x"001a3",
5878=>x"001a3",
5879=>x"001a3",
5880=>x"001a4",
5881=>x"001a4",
5882=>x"001a4",
5883=>x"001a4",
5884=>x"001a4",
5885=>x"001a4",
5886=>x"001a4",
5887=>x"001a4",
5888=>x"001a4",
5889=>x"001a4",
5890=>x"001a4",
5891=>x"001a4",
5892=>x"001a4",
5893=>x"001a4",
5894=>x"001a5",
5895=>x"001a5",
5896=>x"001a5",
5897=>x"001a5",
5898=>x"001a5",
5899=>x"001a5",
5900=>x"001a5",
5901=>x"001a5",
5902=>x"001a5",
5903=>x"001a5",
5904=>x"001a5",
5905=>x"001a5",
5906=>x"001a5",
5907=>x"001a5",
5908=>x"001a6",
5909=>x"001a6",
5910=>x"001a6",
5911=>x"001a6",
5912=>x"001a6",
5913=>x"001a6",
5914=>x"001a6",
5915=>x"001a6",
5916=>x"001a6",
5917=>x"001a6",
5918=>x"001a6",
5919=>x"001a6",
5920=>x"001a6",
5921=>x"001a6",
5922=>x"001a7",
5923=>x"001a7",
5924=>x"001a7",
5925=>x"001a7",
5926=>x"001a7",
5927=>x"001a7",
5928=>x"001a7",
5929=>x"001a7",
5930=>x"001a7",
5931=>x"001a7",
5932=>x"001a7",
5933=>x"001a7",
5934=>x"001a7",
5935=>x"001a7",
5936=>x"001a8",
5937=>x"001a8",
5938=>x"001a8",
5939=>x"001a8",
5940=>x"001a8",
5941=>x"001a8",
5942=>x"001a8",
5943=>x"001a8",
5944=>x"001a8",
5945=>x"001a8",
5946=>x"001a8",
5947=>x"001a8",
5948=>x"001a8",
5949=>x"001a8",
5950=>x"001a9",
5951=>x"001a9",
5952=>x"001a9",
5953=>x"001a9",
5954=>x"001a9",
5955=>x"001a9",
5956=>x"001a9",
5957=>x"001a9",
5958=>x"001a9",
5959=>x"001a9",
5960=>x"001a9",
5961=>x"001a9",
5962=>x"001a9",
5963=>x"001a9",
5964=>x"001aa",
5965=>x"001aa",
5966=>x"001aa",
5967=>x"001aa",
5968=>x"001aa",
5969=>x"001aa",
5970=>x"001aa",
5971=>x"001aa",
5972=>x"001aa",
5973=>x"001aa",
5974=>x"001aa",
5975=>x"001aa",
5976=>x"001aa",
5977=>x"001aa",
5978=>x"001ab",
5979=>x"001ab",
5980=>x"001ab",
5981=>x"001ab",
5982=>x"001ab",
5983=>x"001ab",
5984=>x"001ab",
5985=>x"001ab",
5986=>x"001ab",
5987=>x"001ab",
5988=>x"001ab",
5989=>x"001ab",
5990=>x"001ab",
5991=>x"001ab",
5992=>x"001ac",
5993=>x"001ac",
5994=>x"001ac",
5995=>x"001ac",
5996=>x"001ac",
5997=>x"001ac",
5998=>x"001ac",
5999=>x"001ac",
6000=>x"001ac",
6001=>x"001ac",
6002=>x"001ac",
6003=>x"001ac",
6004=>x"001ac",
6005=>x"001ac",
6006=>x"001ad",
6007=>x"001ad",
6008=>x"001ad",
6009=>x"001ad",
6010=>x"001ad",
6011=>x"001ad",
6012=>x"001ad",
6013=>x"001ad",
6014=>x"001ad",
6015=>x"001ad",
6016=>x"001ad",
6017=>x"001ad",
6018=>x"001ad",
6019=>x"001ad",
6020=>x"001ae",
6021=>x"001ae",
6022=>x"001ae",
6023=>x"001ae",
6024=>x"001ae",
6025=>x"001ae",
6026=>x"001ae",
6027=>x"001ae",
6028=>x"001ae",
6029=>x"001ae",
6030=>x"001ae",
6031=>x"001ae",
6032=>x"001ae",
6033=>x"001ae",
6034=>x"001af",
6035=>x"001af",
6036=>x"001af",
6037=>x"001af",
6038=>x"001af",
6039=>x"001af",
6040=>x"001af",
6041=>x"001af",
6042=>x"001af",
6043=>x"001af",
6044=>x"001af",
6045=>x"001af",
6046=>x"001af",
6047=>x"001af",
6048=>x"001b0",
6049=>x"001b0",
6050=>x"001b0",
6051=>x"001b0",
6052=>x"001b0",
6053=>x"001b0",
6054=>x"001b0",
6055=>x"001b0",
6056=>x"001b0",
6057=>x"001b0",
6058=>x"001b0",
6059=>x"001b0",
6060=>x"001b0",
6061=>x"001b0",
6062=>x"001b1",
6063=>x"001b1",
6064=>x"001b1",
6065=>x"001b1",
6066=>x"001b1",
6067=>x"001b1",
6068=>x"001b1",
6069=>x"001b1",
6070=>x"001b1",
6071=>x"001b1",
6072=>x"001b1",
6073=>x"001b1",
6074=>x"001b1",
6075=>x"001b1",
6076=>x"001b2",
6077=>x"001b2",
6078=>x"001b2",
6079=>x"001b2",
6080=>x"001b2",
6081=>x"001b2",
6082=>x"001b2",
6083=>x"001b2",
6084=>x"001b2",
6085=>x"001b2",
6086=>x"001b2",
6087=>x"001b2",
6088=>x"001b2",
6089=>x"001b2",
6090=>x"001b3",
6091=>x"001b3",
6092=>x"001b3",
6093=>x"001b3",
6094=>x"001b3",
6095=>x"001b3",
6096=>x"001b3",
6097=>x"001b3",
6098=>x"001b3",
6099=>x"001b3",
6100=>x"001b3",
6101=>x"001b3",
6102=>x"001b3",
6103=>x"001b3",
6104=>x"001b4",
6105=>x"001b4",
6106=>x"001b4",
6107=>x"001b4",
6108=>x"001b4",
6109=>x"001b4",
6110=>x"001b4",
6111=>x"001b4",
6112=>x"001b4",
6113=>x"001b4",
6114=>x"001b4",
6115=>x"001b4",
6116=>x"001b4",
6117=>x"001b4",
6118=>x"001b5",
6119=>x"001b5",
6120=>x"001b5",
6121=>x"001b5",
6122=>x"001b5",
6123=>x"001b5",
6124=>x"001b5",
6125=>x"001b5",
6126=>x"001b5",
6127=>x"001b5",
6128=>x"001b5",
6129=>x"001b5",
6130=>x"001b5",
6131=>x"001b5",
6132=>x"001b6",
6133=>x"001b6",
6134=>x"001b6",
6135=>x"001b6",
6136=>x"001b6",
6137=>x"001b6",
6138=>x"001b6",
6139=>x"001b6",
6140=>x"001b6",
6141=>x"001b6",
6142=>x"001b6",
6143=>x"001b6",
6144=>x"001b6",
6145=>x"001b6",
6146=>x"001b7",
6147=>x"001b7",
6148=>x"001b7",
6149=>x"001b7",
6150=>x"001b7",
6151=>x"001b7",
6152=>x"001b7",
6153=>x"001b7",
6154=>x"001b7",
6155=>x"001b7",
6156=>x"001b7",
6157=>x"001b7",
6158=>x"001b7",
6159=>x"001b7",
6160=>x"001b8",
6161=>x"001b8",
6162=>x"001b8",
6163=>x"001b8",
6164=>x"001b8",
6165=>x"001b8",
6166=>x"001b8",
6167=>x"001b8",
6168=>x"001b8",
6169=>x"001b8",
6170=>x"001b8",
6171=>x"001b8",
6172=>x"001b8",
6173=>x"001b8",
6174=>x"001b9",
6175=>x"001b9",
6176=>x"001b9",
6177=>x"001b9",
6178=>x"001b9",
6179=>x"001b9",
6180=>x"001b9",
6181=>x"001b9",
6182=>x"001b9",
6183=>x"001b9",
6184=>x"001b9",
6185=>x"001b9",
6186=>x"001b9",
6187=>x"001b9",
6188=>x"001ba",
6189=>x"001ba",
6190=>x"001ba",
6191=>x"001ba",
6192=>x"001ba",
6193=>x"001ba",
6194=>x"001ba",
6195=>x"001ba",
6196=>x"001ba",
6197=>x"001ba",
6198=>x"001ba",
6199=>x"001ba",
6200=>x"001ba",
6201=>x"001ba",
6202=>x"001bb",
6203=>x"001bb",
6204=>x"001bb",
6205=>x"001bb",
6206=>x"001bb",
6207=>x"001bb",
6208=>x"001bb",
6209=>x"001bb",
6210=>x"001bb",
6211=>x"001bb",
6212=>x"001bb",
6213=>x"001bb",
6214=>x"001bb",
6215=>x"001bb",
6216=>x"001bc",
6217=>x"001bc",
6218=>x"001bc",
6219=>x"001bc",
6220=>x"001bc",
6221=>x"001bc",
6222=>x"001bc",
6223=>x"001bc",
6224=>x"001bc",
6225=>x"001bc",
6226=>x"001bc",
6227=>x"001bc",
6228=>x"001bc",
6229=>x"001bc",
6230=>x"001bd",
6231=>x"001bd",
6232=>x"001bd",
6233=>x"001bd",
6234=>x"001bd",
6235=>x"001bd",
6236=>x"001bd",
6237=>x"001bd",
6238=>x"001bd",
6239=>x"001bd",
6240=>x"001bd",
6241=>x"001bd",
6242=>x"001bd",
6243=>x"001bd",
6244=>x"001be",
6245=>x"001be",
6246=>x"001be",
6247=>x"001be",
6248=>x"001be",
6249=>x"001be",
6250=>x"001be",
6251=>x"001be",
6252=>x"001be",
6253=>x"001be",
6254=>x"001be",
6255=>x"001be",
6256=>x"001be",
6257=>x"001be",
6258=>x"001bf",
6259=>x"001bf",
6260=>x"001bf",
6261=>x"001bf",
6262=>x"001bf",
6263=>x"001bf",
6264=>x"001bf",
6265=>x"001bf",
6266=>x"001bf",
6267=>x"001bf",
6268=>x"001bf",
6269=>x"001bf",
6270=>x"001bf",
6271=>x"001bf",
6272=>x"001c0",
6273=>x"001c0",
6274=>x"001c0",
6275=>x"001c0",
6276=>x"001c0",
6277=>x"001c0",
6278=>x"001c0",
6279=>x"001c0",
6280=>x"001c0",
6281=>x"001c0",
6282=>x"001c0",
6283=>x"001c0",
6284=>x"001c0",
6285=>x"001c0",
6286=>x"001c1",
6287=>x"001c1",
6288=>x"001c1",
6289=>x"001c1",
6290=>x"001c1",
6291=>x"001c1",
6292=>x"001c1",
6293=>x"001c1",
6294=>x"001c1",
6295=>x"001c1",
6296=>x"001c1",
6297=>x"001c1",
6298=>x"001c1",
6299=>x"001c1",
6300=>x"001c2",
6301=>x"001c2",
6302=>x"001c2",
6303=>x"001c2",
6304=>x"001c2",
6305=>x"001c2",
6306=>x"001c2",
6307=>x"001c2",
6308=>x"001c2",
6309=>x"001c2",
6310=>x"001c2",
6311=>x"001c2",
6312=>x"001c2",
6313=>x"001c2",
6314=>x"001c3",
6315=>x"001c3",
6316=>x"001c3",
6317=>x"001c3",
6318=>x"001c3",
6319=>x"001c3",
6320=>x"001c3",
6321=>x"001c3",
6322=>x"001c3",
6323=>x"001c3",
6324=>x"001c3",
6325=>x"001c3",
6326=>x"001c3",
6327=>x"001c3",
6328=>x"001c4",
6329=>x"001c4",
6330=>x"001c4",
6331=>x"001c4",
6332=>x"001c4",
6333=>x"001c4",
6334=>x"001c4",
6335=>x"001c4",
6336=>x"001c4",
6337=>x"001c4",
6338=>x"001c4",
6339=>x"001c4",
6340=>x"001c4",
6341=>x"001c4",
6342=>x"001c5",
6343=>x"001c5",
6344=>x"001c5",
6345=>x"001c5",
6346=>x"001c5",
6347=>x"001c5",
6348=>x"001c5",
6349=>x"001c5",
6350=>x"001c5",
6351=>x"001c5",
6352=>x"001c5",
6353=>x"001c5",
6354=>x"001c5",
6355=>x"001c5",
6356=>x"001c6",
6357=>x"001c6",
6358=>x"001c6",
6359=>x"001c6",
6360=>x"001c6",
6361=>x"001c6",
6362=>x"001c6",
6363=>x"001c6",
6364=>x"001c6",
6365=>x"001c6",
6366=>x"001c6",
6367=>x"001c6",
6368=>x"001c6",
6369=>x"001c6",
6370=>x"001c7",
6371=>x"001c7",
6372=>x"001c7",
6373=>x"001c7",
6374=>x"001c7",
6375=>x"001c7",
6376=>x"001c7",
6377=>x"001c7",
6378=>x"001c7",
6379=>x"001c7",
6380=>x"001c7",
6381=>x"001c7",
6382=>x"001c7",
6383=>x"001c7",
6384=>x"001c8",
6385=>x"001c8",
6386=>x"001c8",
6387=>x"001c8",
6388=>x"001c8",
6389=>x"001c8",
6390=>x"001c8",
6391=>x"001c8",
6392=>x"001c8",
6393=>x"001c8",
6394=>x"001c8",
6395=>x"001c8",
6396=>x"001c8",
6397=>x"001c8",
6398=>x"001c9",
6399=>x"001c9",
6400=>x"001c9",
6401=>x"001c9",
6402=>x"001c9",
6403=>x"001c9",
6404=>x"001c9",
6405=>x"001c9",
6406=>x"001c9",
6407=>x"001c9",
6408=>x"001c9",
6409=>x"001c9",
6410=>x"001c9",
6411=>x"001c9",
6412=>x"001ca",
6413=>x"001ca",
6414=>x"001ca",
6415=>x"001ca",
6416=>x"001ca",
6417=>x"001ca",
6418=>x"001ca",
6419=>x"001ca",
6420=>x"001ca",
6421=>x"001ca",
6422=>x"001ca",
6423=>x"001ca",
6424=>x"001ca",
6425=>x"001ca",
6426=>x"001cb",
6427=>x"001cb",
6428=>x"001cb",
6429=>x"001cb",
6430=>x"001cb",
6431=>x"001cb",
6432=>x"001cb",
6433=>x"001cb",
6434=>x"001cb",
6435=>x"001cb",
6436=>x"001cb",
6437=>x"001cb",
6438=>x"001cb",
6439=>x"001cb",
6440=>x"001cc",
6441=>x"001cc",
6442=>x"001cc",
6443=>x"001cc",
6444=>x"001cc",
6445=>x"001cc",
6446=>x"001cc",
6447=>x"001cc",
6448=>x"001cc",
6449=>x"001cc",
6450=>x"001cc",
6451=>x"001cc",
6452=>x"001cc",
6453=>x"001cc",
6454=>x"001cd",
6455=>x"001cd",
6456=>x"001cd",
6457=>x"001cd",
6458=>x"001cd",
6459=>x"001cd",
6460=>x"001cd",
6461=>x"001cd",
6462=>x"001cd",
6463=>x"001cd",
6464=>x"001cd",
6465=>x"001cd",
6466=>x"001cd",
6467=>x"001cd",
6468=>x"001ce",
6469=>x"001ce",
6470=>x"001ce",
6471=>x"001ce",
6472=>x"001ce",
6473=>x"001ce",
6474=>x"001ce",
6475=>x"001ce",
6476=>x"001ce",
6477=>x"001ce",
6478=>x"001ce",
6479=>x"001ce",
6480=>x"001ce",
6481=>x"001ce",
6482=>x"001cf",
6483=>x"001cf",
6484=>x"001cf",
6485=>x"001cf",
6486=>x"001cf",
6487=>x"001cf",
6488=>x"001cf",
6489=>x"001cf",
6490=>x"001cf",
6491=>x"001cf",
6492=>x"001cf",
6493=>x"001cf",
6494=>x"001cf",
6495=>x"001cf",
6496=>x"001d0",
6497=>x"001d0",
6498=>x"001d0",
6499=>x"001d0",
6500=>x"001d0",
6501=>x"001d0",
6502=>x"001d0",
6503=>x"001d0",
6504=>x"001d0",
6505=>x"001d0",
6506=>x"001d0",
6507=>x"001d0",
6508=>x"001d0",
6509=>x"001d0",
6510=>x"001d1",
6511=>x"001d1",
6512=>x"001d1",
6513=>x"001d1",
6514=>x"001d1",
6515=>x"001d1",
6516=>x"001d1",
6517=>x"001d1",
6518=>x"001d1",
6519=>x"001d1",
6520=>x"001d1",
6521=>x"001d1",
6522=>x"001d1",
6523=>x"001d1",
6524=>x"001d2",
6525=>x"001d2",
6526=>x"001d2",
6527=>x"001d2",
6528=>x"001d2",
6529=>x"001d2",
6530=>x"001d2",
6531=>x"001d2",
6532=>x"001d2",
6533=>x"001d2",
6534=>x"001d2",
6535=>x"001d2",
6536=>x"001d2",
6537=>x"001d2",
6538=>x"001d3",
6539=>x"001d3",
6540=>x"001d3",
6541=>x"001d3",
6542=>x"001d3",
6543=>x"001d3",
6544=>x"001d3",
6545=>x"001d3",
6546=>x"001d3",
6547=>x"001d3",
6548=>x"001d3",
6549=>x"001d3",
6550=>x"001d3",
6551=>x"001d3",
6552=>x"001d4",
6553=>x"001d4",
6554=>x"001d4",
6555=>x"001d4",
6556=>x"001d4",
6557=>x"001d4",
6558=>x"001d4",
6559=>x"001d4",
6560=>x"001d4",
6561=>x"001d4",
6562=>x"001d4",
6563=>x"001d4",
6564=>x"001d4",
6565=>x"001d4",
6566=>x"001d5",
6567=>x"001d5",
6568=>x"001d5",
6569=>x"001d5",
6570=>x"001d5",
6571=>x"001d5",
6572=>x"001d5",
6573=>x"001d5",
6574=>x"001d5",
6575=>x"001d5",
6576=>x"001d5",
6577=>x"001d5",
6578=>x"001d5",
6579=>x"001d5",
6580=>x"001d6",
6581=>x"001d6",
6582=>x"001d6",
6583=>x"001d6",
6584=>x"001d6",
6585=>x"001d6",
6586=>x"001d6",
6587=>x"001d6",
6588=>x"001d6",
6589=>x"001d6",
6590=>x"001d6",
6591=>x"001d6",
6592=>x"001d6",
6593=>x"001d6",
6594=>x"001d7",
6595=>x"001d7",
6596=>x"001d7",
6597=>x"001d7",
6598=>x"001d7",
6599=>x"001d7",
6600=>x"001d7",
6601=>x"001d7",
6602=>x"001d7",
6603=>x"001d7",
6604=>x"001d7",
6605=>x"001d7",
6606=>x"001d7",
6607=>x"001d7",
6608=>x"001d8",
6609=>x"001d8",
6610=>x"001d8",
6611=>x"001d8",
6612=>x"001d8",
6613=>x"001d8",
6614=>x"001d8",
6615=>x"001d8",
6616=>x"001d8",
6617=>x"001d8",
6618=>x"001d8",
6619=>x"001d8",
6620=>x"001d8",
6621=>x"001d8",
6622=>x"001d9",
6623=>x"001d9",
6624=>x"001d9",
6625=>x"001d9",
6626=>x"001d9",
6627=>x"001d9",
6628=>x"001d9",
6629=>x"001d9",
6630=>x"001d9",
6631=>x"001d9",
6632=>x"001d9",
6633=>x"001d9",
6634=>x"001d9",
6635=>x"001d9",
6636=>x"001da",
6637=>x"001da",
6638=>x"001da",
6639=>x"001da",
6640=>x"001da",
6641=>x"001da",
6642=>x"001da",
6643=>x"001da",
6644=>x"001da",
6645=>x"001da",
6646=>x"001da",
6647=>x"001da",
6648=>x"001da",
6649=>x"001da",
6650=>x"001db",
6651=>x"001db",
6652=>x"001db",
6653=>x"001db",
6654=>x"001db",
6655=>x"001db",
6656=>x"001db",
6657=>x"001db",
6658=>x"001db",
6659=>x"001db",
6660=>x"001db",
6661=>x"001db",
6662=>x"001db",
6663=>x"001db",
6664=>x"001dc",
6665=>x"001dc",
6666=>x"001dc",
6667=>x"001dc",
6668=>x"001dc",
6669=>x"001dc",
6670=>x"001dc",
6671=>x"001dc",
6672=>x"001dc",
6673=>x"001dc",
6674=>x"001dc",
6675=>x"001dc",
6676=>x"001dc",
6677=>x"001dc",
6678=>x"001dd",
6679=>x"001dd",
6680=>x"001dd",
6681=>x"001dd",
6682=>x"001dd",
6683=>x"001dd",
6684=>x"001dd",
6685=>x"001dd",
6686=>x"001dd",
6687=>x"001dd",
6688=>x"001dd",
6689=>x"001dd",
6690=>x"001dd",
6691=>x"001dd",
6692=>x"001de",
6693=>x"001de",
6694=>x"001de",
6695=>x"001de",
6696=>x"001de",
6697=>x"001de",
6698=>x"001de",
6699=>x"001de",
6700=>x"001de",
6701=>x"001de",
6702=>x"001de",
6703=>x"001de",
6704=>x"001de",
6705=>x"001de",
6706=>x"001df",
6707=>x"001df",
6708=>x"001df",
6709=>x"001df",
6710=>x"001df",
6711=>x"001df",
6712=>x"001df",
6713=>x"001df",
6714=>x"001df",
6715=>x"001df",
6716=>x"001df",
6717=>x"001df",
6718=>x"001df",
6719=>x"001df",
6720=>x"001e0",
6721=>x"001e0",
6722=>x"001e0",
6723=>x"001e0",
6724=>x"001e0",
6725=>x"001e0",
6726=>x"001e0",
6727=>x"001e0",
6728=>x"001e0",
6729=>x"001e0",
6730=>x"001e0",
6731=>x"001e0",
6732=>x"001e0",
6733=>x"001e0",
6734=>x"001e1",
6735=>x"001e1",
6736=>x"001e1",
6737=>x"001e1",
6738=>x"001e1",
6739=>x"001e1",
6740=>x"001e1",
6741=>x"001e1",
6742=>x"001e1",
6743=>x"001e1",
6744=>x"001e1",
6745=>x"001e1",
6746=>x"001e1",
6747=>x"001e1",
6748=>x"001e2",
6749=>x"001e2",
6750=>x"001e2",
6751=>x"001e2",
6752=>x"001e2",
6753=>x"001e2",
6754=>x"001e2",
6755=>x"001e2",
6756=>x"001e2",
6757=>x"001e2",
6758=>x"001e2",
6759=>x"001e2",
6760=>x"001e2",
6761=>x"001e2",
6762=>x"001e3",
6763=>x"001e3",
6764=>x"001e3",
6765=>x"001e3",
6766=>x"001e3",
6767=>x"001e3",
6768=>x"001e3",
6769=>x"001e3",
6770=>x"001e3",
6771=>x"001e3",
6772=>x"001e3",
6773=>x"001e3",
6774=>x"001e3",
6775=>x"001e3",
6776=>x"001e4",
6777=>x"001e4",
6778=>x"001e4",
6779=>x"001e4",
6780=>x"001e4",
6781=>x"001e4",
6782=>x"001e4",
6783=>x"001e4",
6784=>x"001e4",
6785=>x"001e4",
6786=>x"001e4",
6787=>x"001e4",
6788=>x"001e4",
6789=>x"001e4",
6790=>x"001e5",
6791=>x"001e5",
6792=>x"001e5",
6793=>x"001e5",
6794=>x"001e5",
6795=>x"001e5",
6796=>x"001e5",
6797=>x"001e5",
6798=>x"001e5",
6799=>x"001e5",
6800=>x"001e5",
6801=>x"001e5",
6802=>x"001e5",
6803=>x"001e5",
6804=>x"001e6",
6805=>x"001e6",
6806=>x"001e6",
6807=>x"001e6",
6808=>x"001e6",
6809=>x"001e6",
6810=>x"001e6",
6811=>x"001e6",
6812=>x"001e6",
6813=>x"001e6",
6814=>x"001e6",
6815=>x"001e6",
6816=>x"001e6",
6817=>x"001e6",
6818=>x"001e7",
6819=>x"001e7",
6820=>x"001e7",
6821=>x"001e7",
6822=>x"001e7",
6823=>x"001e7",
6824=>x"001e7",
6825=>x"001e7",
6826=>x"001e7",
6827=>x"001e7",
6828=>x"001e7",
6829=>x"001e7",
6830=>x"001e7",
6831=>x"001e7",
6832=>x"001e8",
6833=>x"001e8",
6834=>x"001e8",
6835=>x"001e8",
6836=>x"001e8",
6837=>x"001e8",
6838=>x"001e8",
6839=>x"001e8",
6840=>x"001e8",
6841=>x"001e8",
6842=>x"001e8",
6843=>x"001e8",
6844=>x"001e8",
6845=>x"001e8",
6846=>x"001e9",
6847=>x"001e9",
6848=>x"001e9",
6849=>x"001e9",
6850=>x"001e9",
6851=>x"001e9",
6852=>x"001e9",
6853=>x"001e9",
6854=>x"001e9",
6855=>x"001e9",
6856=>x"001e9",
6857=>x"001e9",
6858=>x"001e9",
6859=>x"001e9",
6860=>x"001ea",
6861=>x"001ea",
6862=>x"001ea",
6863=>x"001ea",
6864=>x"001ea",
6865=>x"001ea",
6866=>x"001ea",
6867=>x"001ea",
6868=>x"001ea",
6869=>x"001ea",
6870=>x"001ea",
6871=>x"001ea",
6872=>x"001ea",
6873=>x"001ea",
6874=>x"001eb",
6875=>x"001eb",
6876=>x"001eb",
6877=>x"001eb",
6878=>x"001eb",
6879=>x"001eb",
6880=>x"001eb",
6881=>x"001eb",
6882=>x"001eb",
6883=>x"001eb",
6884=>x"001eb",
6885=>x"001eb",
6886=>x"001eb",
6887=>x"001eb",
6888=>x"001ec",
6889=>x"001ec",
6890=>x"001ec",
6891=>x"001ec",
6892=>x"001ec",
6893=>x"001ec",
6894=>x"001ec",
6895=>x"001ec",
6896=>x"001ec",
6897=>x"001ec",
6898=>x"001ec",
6899=>x"001ec",
6900=>x"001ec",
6901=>x"001ec",
6902=>x"001ed",
6903=>x"001ed",
6904=>x"001ed",
6905=>x"001ed",
6906=>x"001ed",
6907=>x"001ed",
6908=>x"001ed",
6909=>x"001ed",
6910=>x"001ed",
6911=>x"001ed",
6912=>x"001ed",
6913=>x"001ed",
6914=>x"001ed",
6915=>x"001ed",
6916=>x"001ee",
6917=>x"001ee",
6918=>x"001ee",
6919=>x"001ee",
6920=>x"001ee",
6921=>x"001ee",
6922=>x"001ee",
6923=>x"001ee",
6924=>x"001ee",
6925=>x"001ee",
6926=>x"001ee",
6927=>x"001ee",
6928=>x"001ee",
6929=>x"001ee",
6930=>x"001ef",
6931=>x"001ef",
6932=>x"001ef",
6933=>x"001ef",
6934=>x"001ef",
6935=>x"001ef",
6936=>x"001ef",
6937=>x"001ef",
6938=>x"001ef",
6939=>x"001ef",
6940=>x"001ef",
6941=>x"001ef",
6942=>x"001ef",
6943=>x"001ef",
6944=>x"001f0",
6945=>x"001f0",
6946=>x"001f0",
6947=>x"001f0",
6948=>x"001f0",
6949=>x"001f0",
6950=>x"001f0",
6951=>x"001f0",
6952=>x"001f0",
6953=>x"001f0",
6954=>x"001f0",
6955=>x"001f0",
6956=>x"001f0",
6957=>x"001f0",
6958=>x"001f1",
6959=>x"001f1",
6960=>x"001f1",
6961=>x"001f1",
6962=>x"001f1",
6963=>x"001f1",
6964=>x"001f1",
6965=>x"001f1",
6966=>x"001f1",
6967=>x"001f1",
6968=>x"001f1",
6969=>x"001f1",
6970=>x"001f1",
6971=>x"001f1",
6972=>x"001f2",
6973=>x"001f2",
6974=>x"001f2",
6975=>x"001f2",
6976=>x"001f2",
6977=>x"001f2",
6978=>x"001f2",
6979=>x"001f2",
6980=>x"001f2",
6981=>x"001f2",
6982=>x"001f2",
6983=>x"001f2",
6984=>x"001f2",
6985=>x"001f2",
6986=>x"001f3",
6987=>x"001f3",
6988=>x"001f3",
6989=>x"001f3",
6990=>x"001f3",
6991=>x"001f3",
6992=>x"001f3",
6993=>x"001f3",
6994=>x"001f3",
6995=>x"001f3",
6996=>x"001f3",
6997=>x"001f3",
6998=>x"001f3",
6999=>x"001f3",
7000=>x"001f4",
7001=>x"001f4",
7002=>x"001f4",
7003=>x"001f4",
7004=>x"001f4",
7005=>x"001f4",
7006=>x"001f4",
7007=>x"001f4",
7008=>x"001f4",
7009=>x"001f4",
7010=>x"001f4",
7011=>x"001f4",
7012=>x"001f4",
7013=>x"001f4",
7014=>x"001f5",
7015=>x"001f5",
7016=>x"001f5",
7017=>x"001f5",
7018=>x"001f5",
7019=>x"001f5",
7020=>x"001f5",
7021=>x"001f5",
7022=>x"001f5",
7023=>x"001f5",
7024=>x"001f5",
7025=>x"001f5",
7026=>x"001f5",
7027=>x"001f5",
7028=>x"001f6",
7029=>x"001f6",
7030=>x"001f6",
7031=>x"001f6",
7032=>x"001f6",
7033=>x"001f6",
7034=>x"001f6",
7035=>x"001f6",
7036=>x"001f6",
7037=>x"001f6",
7038=>x"001f6",
7039=>x"001f6",
7040=>x"001f6",
7041=>x"001f6",
7042=>x"001f7",
7043=>x"001f7",
7044=>x"001f7",
7045=>x"001f7",
7046=>x"001f7",
7047=>x"001f7",
7048=>x"001f7",
7049=>x"001f7",
7050=>x"001f7",
7051=>x"001f7",
7052=>x"001f7",
7053=>x"001f7",
7054=>x"001f7",
7055=>x"001f7",
7056=>x"001f8",
7057=>x"001f8",
7058=>x"001f8",
7059=>x"001f8",
7060=>x"001f8",
7061=>x"001f8",
7062=>x"001f8",
7063=>x"001f8",
7064=>x"001f8",
7065=>x"001f8",
7066=>x"001f8",
7067=>x"001f8",
7068=>x"001f8",
7069=>x"001f8",
7070=>x"001f9",
7071=>x"001f9",
7072=>x"001f9",
7073=>x"001f9",
7074=>x"001f9",
7075=>x"001f9",
7076=>x"001f9",
7077=>x"001f9",
7078=>x"001f9",
7079=>x"001f9",
7080=>x"001f9",
7081=>x"001f9",
7082=>x"001f9",
7083=>x"001f9",
7084=>x"001fa",
7085=>x"001fa",
7086=>x"001fa",
7087=>x"001fa",
7088=>x"001fa",
7089=>x"001fa",
7090=>x"001fa",
7091=>x"001fa",
7092=>x"001fa",
7093=>x"001fa",
7094=>x"001fa",
7095=>x"001fa",
7096=>x"001fa",
7097=>x"001fa",
7098=>x"001fb",
7099=>x"001fb",
7100=>x"001fb",
7101=>x"001fb",
7102=>x"001fb",
7103=>x"001fb",
7104=>x"001fb",
7105=>x"001fb",
7106=>x"001fb",
7107=>x"001fb",
7108=>x"001fb",
7109=>x"001fb",
7110=>x"001fb",
7111=>x"001fb",
7112=>x"001fc",
7113=>x"001fc",
7114=>x"001fc",
7115=>x"001fc",
7116=>x"001fc",
7117=>x"001fc",
7118=>x"001fc",
7119=>x"001fc",
7120=>x"001fc",
7121=>x"001fc",
7122=>x"001fc",
7123=>x"001fc",
7124=>x"001fc",
7125=>x"001fc",
7126=>x"001fd",
7127=>x"001fd",
7128=>x"001fd",
7129=>x"001fd",
7130=>x"001fd",
7131=>x"001fd",
7132=>x"001fd",
7133=>x"001fd",
7134=>x"001fd",
7135=>x"001fd",
7136=>x"001fd",
7137=>x"001fd",
7138=>x"001fd",
7139=>x"001fd",
7140=>x"001fe",
7141=>x"001fe",
7142=>x"001fe",
7143=>x"001fe",
7144=>x"001fe",
7145=>x"001fe",
7146=>x"001fe",
7147=>x"001fe",
7148=>x"001fe",
7149=>x"001fe",
7150=>x"001fe",
7151=>x"001fe",
7152=>x"001fe",
7153=>x"001fe",
7154=>x"001ff",
7155=>x"001ff",
7156=>x"001ff",
7157=>x"001ff",
7158=>x"001ff",
7159=>x"001ff",
7160=>x"001ff",
7161=>x"001ff",
7162=>x"001ff",
7163=>x"001ff",
7164=>x"001ff",
7165=>x"001ff",
7166=>x"001ff",
7167=>x"001ff",
7168=>x"00200",
7169=>x"00200",
7170=>x"00200",
7171=>x"00200",
7172=>x"00200",
7173=>x"00200",
7174=>x"00200",
7175=>x"00200",
7176=>x"00200",
7177=>x"00200",
7178=>x"00200",
7179=>x"00200",
7180=>x"00200",
7181=>x"00200",
7182=>x"00201",
7183=>x"00201",
7184=>x"00201",
7185=>x"00201",
7186=>x"00201",
7187=>x"00201",
7188=>x"00201",
7189=>x"00201",
7190=>x"00201",
7191=>x"00201",
7192=>x"00201",
7193=>x"00201",
7194=>x"00201",
7195=>x"00201",
7196=>x"00202",
7197=>x"00202",
7198=>x"00202",
7199=>x"00202",
7200=>x"00202",
7201=>x"00202",
7202=>x"00202",
7203=>x"00202",
7204=>x"00202",
7205=>x"00202",
7206=>x"00202",
7207=>x"00202",
7208=>x"00202",
7209=>x"00202",
7210=>x"00203",
7211=>x"00203",
7212=>x"00203",
7213=>x"00203",
7214=>x"00203",
7215=>x"00203",
7216=>x"00203",
7217=>x"00203",
7218=>x"00203",
7219=>x"00203",
7220=>x"00203",
7221=>x"00203",
7222=>x"00203",
7223=>x"00203",
7224=>x"00204",
7225=>x"00204",
7226=>x"00204",
7227=>x"00204",
7228=>x"00204",
7229=>x"00204",
7230=>x"00204",
7231=>x"00204",
7232=>x"00204",
7233=>x"00204",
7234=>x"00204",
7235=>x"00204",
7236=>x"00204",
7237=>x"00204",
7238=>x"00205",
7239=>x"00205",
7240=>x"00205",
7241=>x"00205",
7242=>x"00205",
7243=>x"00205",
7244=>x"00205",
7245=>x"00205",
7246=>x"00205",
7247=>x"00205",
7248=>x"00205",
7249=>x"00205",
7250=>x"00205",
7251=>x"00205",
7252=>x"00206",
7253=>x"00206",
7254=>x"00206",
7255=>x"00206",
7256=>x"00206",
7257=>x"00206",
7258=>x"00206",
7259=>x"00206",
7260=>x"00206",
7261=>x"00206",
7262=>x"00206",
7263=>x"00206",
7264=>x"00206",
7265=>x"00206",
7266=>x"00207",
7267=>x"00207",
7268=>x"00207",
7269=>x"00207",
7270=>x"00207",
7271=>x"00207",
7272=>x"00207",
7273=>x"00207",
7274=>x"00207",
7275=>x"00207",
7276=>x"00207",
7277=>x"00207",
7278=>x"00207",
7279=>x"00207",
7280=>x"00208",
7281=>x"00208",
7282=>x"00208",
7283=>x"00208",
7284=>x"00208",
7285=>x"00208",
7286=>x"00208",
7287=>x"00208",
7288=>x"00208",
7289=>x"00208",
7290=>x"00208",
7291=>x"00208",
7292=>x"00208",
7293=>x"00208",
7294=>x"00209",
7295=>x"00209",
7296=>x"00209",
7297=>x"00209",
7298=>x"00209",
7299=>x"00209",
7300=>x"00209",
7301=>x"00209",
7302=>x"00209",
7303=>x"00209",
7304=>x"00209",
7305=>x"00209",
7306=>x"00209",
7307=>x"00209",
7308=>x"0020a",
7309=>x"0020a",
7310=>x"0020a",
7311=>x"0020a",
7312=>x"0020a",
7313=>x"0020a",
7314=>x"0020a",
7315=>x"0020a",
7316=>x"0020a",
7317=>x"0020a",
7318=>x"0020a",
7319=>x"0020a",
7320=>x"0020a",
7321=>x"0020a",
7322=>x"0020b",
7323=>x"0020b",
7324=>x"0020b",
7325=>x"0020b",
7326=>x"0020b",
7327=>x"0020b",
7328=>x"0020b",
7329=>x"0020b",
7330=>x"0020b",
7331=>x"0020b",
7332=>x"0020b",
7333=>x"0020b",
7334=>x"0020b",
7335=>x"0020b",
7336=>x"0020c",
7337=>x"0020c",
7338=>x"0020c",
7339=>x"0020c",
7340=>x"0020c",
7341=>x"0020c",
7342=>x"0020c",
7343=>x"0020c",
7344=>x"0020c",
7345=>x"0020c",
7346=>x"0020c",
7347=>x"0020c",
7348=>x"0020c",
7349=>x"0020c",
7350=>x"0020d",
7351=>x"0020d",
7352=>x"0020d",
7353=>x"0020d",
7354=>x"0020d",
7355=>x"0020d",
7356=>x"0020d",
7357=>x"0020d",
7358=>x"0020d",
7359=>x"0020d",
7360=>x"0020d",
7361=>x"0020d",
7362=>x"0020d",
7363=>x"0020d",
7364=>x"0020e",
7365=>x"0020e",
7366=>x"0020e",
7367=>x"0020e",
7368=>x"0020e",
7369=>x"0020e",
7370=>x"0020e",
7371=>x"0020e",
7372=>x"0020e",
7373=>x"0020e",
7374=>x"0020e",
7375=>x"0020e",
7376=>x"0020e",
7377=>x"0020e",
7378=>x"0020f",
7379=>x"0020f",
7380=>x"0020f",
7381=>x"0020f",
7382=>x"0020f",
7383=>x"0020f",
7384=>x"0020f",
7385=>x"0020f",
7386=>x"0020f",
7387=>x"0020f",
7388=>x"0020f",
7389=>x"0020f",
7390=>x"0020f",
7391=>x"0020f",
7392=>x"00210",
7393=>x"00210",
7394=>x"00210",
7395=>x"00210",
7396=>x"00210",
7397=>x"00210",
7398=>x"00210",
7399=>x"00210",
7400=>x"00210",
7401=>x"00210",
7402=>x"00210",
7403=>x"00210",
7404=>x"00210",
7405=>x"00210",
7406=>x"00211",
7407=>x"00211",
7408=>x"00211",
7409=>x"00211",
7410=>x"00211",
7411=>x"00211",
7412=>x"00211",
7413=>x"00211",
7414=>x"00211",
7415=>x"00211",
7416=>x"00211",
7417=>x"00211",
7418=>x"00211",
7419=>x"00211",
7420=>x"00212",
7421=>x"00212",
7422=>x"00212",
7423=>x"00212",
7424=>x"00212",
7425=>x"00212",
7426=>x"00212",
7427=>x"00212",
7428=>x"00212",
7429=>x"00212",
7430=>x"00212",
7431=>x"00212",
7432=>x"00212",
7433=>x"00212",
7434=>x"00213",
7435=>x"00213",
7436=>x"00213",
7437=>x"00213",
7438=>x"00213",
7439=>x"00213",
7440=>x"00213",
7441=>x"00213",
7442=>x"00213",
7443=>x"00213",
7444=>x"00213",
7445=>x"00213",
7446=>x"00213",
7447=>x"00213",
7448=>x"00214",
7449=>x"00214",
7450=>x"00214",
7451=>x"00214",
7452=>x"00214",
7453=>x"00214",
7454=>x"00214",
7455=>x"00214",
7456=>x"00214",
7457=>x"00214",
7458=>x"00214",
7459=>x"00214",
7460=>x"00214",
7461=>x"00214",
7462=>x"00215",
7463=>x"00215",
7464=>x"00215",
7465=>x"00215",
7466=>x"00215",
7467=>x"00215",
7468=>x"00215",
7469=>x"00215",
7470=>x"00215",
7471=>x"00215",
7472=>x"00215",
7473=>x"00215",
7474=>x"00215",
7475=>x"00215",
7476=>x"00216",
7477=>x"00216",
7478=>x"00216",
7479=>x"00216",
7480=>x"00216",
7481=>x"00216",
7482=>x"00216",
7483=>x"00216",
7484=>x"00216",
7485=>x"00216",
7486=>x"00216",
7487=>x"00216",
7488=>x"00216",
7489=>x"00216",
7490=>x"00217",
7491=>x"00217",
7492=>x"00217",
7493=>x"00217",
7494=>x"00217",
7495=>x"00217",
7496=>x"00217",
7497=>x"00217",
7498=>x"00217",
7499=>x"00217",
7500=>x"00217",
7501=>x"00217",
7502=>x"00217",
7503=>x"00217",
7504=>x"00218",
7505=>x"00218",
7506=>x"00218",
7507=>x"00218",
7508=>x"00218",
7509=>x"00218",
7510=>x"00218",
7511=>x"00218",
7512=>x"00218",
7513=>x"00218",
7514=>x"00218",
7515=>x"00218",
7516=>x"00218",
7517=>x"00218",
7518=>x"00219",
7519=>x"00219",
7520=>x"00219",
7521=>x"00219",
7522=>x"00219",
7523=>x"00219",
7524=>x"00219",
7525=>x"00219",
7526=>x"00219",
7527=>x"00219",
7528=>x"00219",
7529=>x"00219",
7530=>x"00219",
7531=>x"00219",
7532=>x"0021a",
7533=>x"0021a",
7534=>x"0021a",
7535=>x"0021a",
7536=>x"0021a",
7537=>x"0021a",
7538=>x"0021a",
7539=>x"0021a",
7540=>x"0021a",
7541=>x"0021a",
7542=>x"0021a",
7543=>x"0021a",
7544=>x"0021a",
7545=>x"0021a",
7546=>x"0021b",
7547=>x"0021b",
7548=>x"0021b",
7549=>x"0021b",
7550=>x"0021b",
7551=>x"0021b",
7552=>x"0021b",
7553=>x"0021b",
7554=>x"0021b",
7555=>x"0021b",
7556=>x"0021b",
7557=>x"0021b",
7558=>x"0021b",
7559=>x"0021b",
7560=>x"0021c",
7561=>x"0021c",
7562=>x"0021c",
7563=>x"0021c",
7564=>x"0021c",
7565=>x"0021c",
7566=>x"0021c",
7567=>x"0021c",
7568=>x"0021c",
7569=>x"0021c",
7570=>x"0021c",
7571=>x"0021c",
7572=>x"0021c",
7573=>x"0021c",
7574=>x"0021d",
7575=>x"0021d",
7576=>x"0021d",
7577=>x"0021d",
7578=>x"0021d",
7579=>x"0021d",
7580=>x"0021d",
7581=>x"0021d",
7582=>x"0021d",
7583=>x"0021d",
7584=>x"0021d",
7585=>x"0021d",
7586=>x"0021d",
7587=>x"0021d",
7588=>x"0021e",
7589=>x"0021e",
7590=>x"0021e",
7591=>x"0021e",
7592=>x"0021e",
7593=>x"0021e",
7594=>x"0021e",
7595=>x"0021e",
7596=>x"0021e",
7597=>x"0021e",
7598=>x"0021e",
7599=>x"0021e",
7600=>x"0021e",
7601=>x"0021e",
7602=>x"0021f",
7603=>x"0021f",
7604=>x"0021f",
7605=>x"0021f",
7606=>x"0021f",
7607=>x"0021f",
7608=>x"0021f",
7609=>x"0021f",
7610=>x"0021f",
7611=>x"0021f",
7612=>x"0021f",
7613=>x"0021f",
7614=>x"0021f",
7615=>x"0021f",
7616=>x"00220",
7617=>x"00220",
7618=>x"00220",
7619=>x"00220",
7620=>x"00220",
7621=>x"00220",
7622=>x"00220",
7623=>x"00220",
7624=>x"00220",
7625=>x"00220",
7626=>x"00220",
7627=>x"00220",
7628=>x"00220",
7629=>x"00220",
7630=>x"00221",
7631=>x"00221",
7632=>x"00221",
7633=>x"00221",
7634=>x"00221",
7635=>x"00221",
7636=>x"00221",
7637=>x"00221",
7638=>x"00221",
7639=>x"00221",
7640=>x"00221",
7641=>x"00221",
7642=>x"00221",
7643=>x"00221",
7644=>x"00222",
7645=>x"00222",
7646=>x"00222",
7647=>x"00222",
7648=>x"00222",
7649=>x"00222",
7650=>x"00222",
7651=>x"00222",
7652=>x"00222",
7653=>x"00222",
7654=>x"00222",
7655=>x"00222",
7656=>x"00222",
7657=>x"00222",
7658=>x"00223",
7659=>x"00223",
7660=>x"00223",
7661=>x"00223",
7662=>x"00223",
7663=>x"00223",
7664=>x"00223",
7665=>x"00223",
7666=>x"00223",
7667=>x"00223",
7668=>x"00223",
7669=>x"00223",
7670=>x"00223",
7671=>x"00223",
7672=>x"00224",
7673=>x"00224",
7674=>x"00224",
7675=>x"00224",
7676=>x"00224",
7677=>x"00224",
7678=>x"00224",
7679=>x"00224",
7680=>x"00224",
7681=>x"00224",
7682=>x"00224",
7683=>x"00224",
7684=>x"00224",
7685=>x"00224",
7686=>x"00225",
7687=>x"00225",
7688=>x"00225",
7689=>x"00225",
7690=>x"00225",
7691=>x"00225",
7692=>x"00225",
7693=>x"00225",
7694=>x"00225",
7695=>x"00225",
7696=>x"00225",
7697=>x"00225",
7698=>x"00225",
7699=>x"00225",
7700=>x"00226",
7701=>x"00226",
7702=>x"00226",
7703=>x"00226",
7704=>x"00226",
7705=>x"00226",
7706=>x"00226",
7707=>x"00226",
7708=>x"00226",
7709=>x"00226",
7710=>x"00226",
7711=>x"00226",
7712=>x"00226",
7713=>x"00226",
7714=>x"00227",
7715=>x"00227",
7716=>x"00227",
7717=>x"00227",
7718=>x"00227",
7719=>x"00227",
7720=>x"00227",
7721=>x"00227",
7722=>x"00227",
7723=>x"00227",
7724=>x"00227",
7725=>x"00227",
7726=>x"00227",
7727=>x"00227",
7728=>x"00228",
7729=>x"00228",
7730=>x"00228",
7731=>x"00228",
7732=>x"00228",
7733=>x"00228",
7734=>x"00228",
7735=>x"00228",
7736=>x"00228",
7737=>x"00228",
7738=>x"00228",
7739=>x"00228",
7740=>x"00228",
7741=>x"00228",
7742=>x"00229",
7743=>x"00229",
7744=>x"00229",
7745=>x"00229",
7746=>x"00229",
7747=>x"00229",
7748=>x"00229",
7749=>x"00229",
7750=>x"00229",
7751=>x"00229",
7752=>x"00229",
7753=>x"00229",
7754=>x"00229",
7755=>x"00229",
7756=>x"0022a",
7757=>x"0022a",
7758=>x"0022a",
7759=>x"0022a",
7760=>x"0022a",
7761=>x"0022a",
7762=>x"0022a",
7763=>x"0022a",
7764=>x"0022a",
7765=>x"0022a",
7766=>x"0022a",
7767=>x"0022a",
7768=>x"0022a",
7769=>x"0022a",
7770=>x"0022b",
7771=>x"0022b",
7772=>x"0022b",
7773=>x"0022b",
7774=>x"0022b",
7775=>x"0022b",
7776=>x"0022b",
7777=>x"0022b",
7778=>x"0022b",
7779=>x"0022b",
7780=>x"0022b",
7781=>x"0022b",
7782=>x"0022b",
7783=>x"0022b",
7784=>x"0022c",
7785=>x"0022c",
7786=>x"0022c",
7787=>x"0022c",
7788=>x"0022c",
7789=>x"0022c",
7790=>x"0022c",
7791=>x"0022c",
7792=>x"0022c",
7793=>x"0022c",
7794=>x"0022c",
7795=>x"0022c",
7796=>x"0022c",
7797=>x"0022c",
7798=>x"0022d",
7799=>x"0022d",
7800=>x"0022d",
7801=>x"0022d",
7802=>x"0022d",
7803=>x"0022d",
7804=>x"0022d",
7805=>x"0022d",
7806=>x"0022d",
7807=>x"0022d",
7808=>x"0022d",
7809=>x"0022d",
7810=>x"0022d",
7811=>x"0022d",
7812=>x"0022e",
7813=>x"0022e",
7814=>x"0022e",
7815=>x"0022e",
7816=>x"0022e",
7817=>x"0022e",
7818=>x"0022e",
7819=>x"0022e",
7820=>x"0022e",
7821=>x"0022e",
7822=>x"0022e",
7823=>x"0022e",
7824=>x"0022e",
7825=>x"0022e",
7826=>x"0022f",
7827=>x"0022f",
7828=>x"0022f",
7829=>x"0022f",
7830=>x"0022f",
7831=>x"0022f",
7832=>x"0022f",
7833=>x"0022f",
7834=>x"0022f",
7835=>x"0022f",
7836=>x"0022f",
7837=>x"0022f",
7838=>x"0022f",
7839=>x"0022f",
7840=>x"00230",
7841=>x"00230",
7842=>x"00230",
7843=>x"00230",
7844=>x"00230",
7845=>x"00230",
7846=>x"00230",
7847=>x"00230",
7848=>x"00230",
7849=>x"00230",
7850=>x"00230",
7851=>x"00230",
7852=>x"00230",
7853=>x"00230",
7854=>x"00231",
7855=>x"00231",
7856=>x"00231",
7857=>x"00231",
7858=>x"00231",
7859=>x"00231",
7860=>x"00231",
7861=>x"00231",
7862=>x"00231",
7863=>x"00231",
7864=>x"00231",
7865=>x"00231",
7866=>x"00231",
7867=>x"00231",
7868=>x"00232",
7869=>x"00232",
7870=>x"00232",
7871=>x"00232",
7872=>x"00232",
7873=>x"00232",
7874=>x"00232",
7875=>x"00232",
7876=>x"00232",
7877=>x"00232",
7878=>x"00232",
7879=>x"00232",
7880=>x"00232",
7881=>x"00232",
7882=>x"00233",
7883=>x"00233",
7884=>x"00233",
7885=>x"00233",
7886=>x"00233",
7887=>x"00233",
7888=>x"00233",
7889=>x"00233",
7890=>x"00233",
7891=>x"00233",
7892=>x"00233",
7893=>x"00233",
7894=>x"00233",
7895=>x"00233",
7896=>x"00234",
7897=>x"00234",
7898=>x"00234",
7899=>x"00234",
7900=>x"00234",
7901=>x"00234",
7902=>x"00234",
7903=>x"00234",
7904=>x"00234",
7905=>x"00234",
7906=>x"00234",
7907=>x"00234",
7908=>x"00234",
7909=>x"00234",
7910=>x"00235",
7911=>x"00235",
7912=>x"00235",
7913=>x"00235",
7914=>x"00235",
7915=>x"00235",
7916=>x"00235",
7917=>x"00235",
7918=>x"00235",
7919=>x"00235",
7920=>x"00235",
7921=>x"00235",
7922=>x"00235",
7923=>x"00235",
7924=>x"00236",
7925=>x"00236",
7926=>x"00236",
7927=>x"00236",
7928=>x"00236",
7929=>x"00236",
7930=>x"00236",
7931=>x"00236",
7932=>x"00236",
7933=>x"00236",
7934=>x"00236",
7935=>x"00236",
7936=>x"00236",
7937=>x"00236",
7938=>x"00237",
7939=>x"00237",
7940=>x"00237",
7941=>x"00237",
7942=>x"00237",
7943=>x"00237",
7944=>x"00237",
7945=>x"00237",
7946=>x"00237",
7947=>x"00237",
7948=>x"00237",
7949=>x"00237",
7950=>x"00237",
7951=>x"00237",
7952=>x"00238",
7953=>x"00238",
7954=>x"00238",
7955=>x"00238",
7956=>x"00238",
7957=>x"00238",
7958=>x"00238",
7959=>x"00238",
7960=>x"00238",
7961=>x"00238",
7962=>x"00238",
7963=>x"00238",
7964=>x"00238",
7965=>x"00238",
7966=>x"00239",
7967=>x"00239",
7968=>x"00239",
7969=>x"00239",
7970=>x"00239",
7971=>x"00239",
7972=>x"00239",
7973=>x"00239",
7974=>x"00239",
7975=>x"00239",
7976=>x"00239",
7977=>x"00239",
7978=>x"00239",
7979=>x"00239",
7980=>x"0023a",
7981=>x"0023a",
7982=>x"0023a",
7983=>x"0023a",
7984=>x"0023a",
7985=>x"0023a",
7986=>x"0023a",
7987=>x"0023a",
7988=>x"0023a",
7989=>x"0023a",
7990=>x"0023a",
7991=>x"0023a",
7992=>x"0023a",
7993=>x"0023a",
7994=>x"0023b",
7995=>x"0023b",
7996=>x"0023b",
7997=>x"0023b",
7998=>x"0023b",
7999=>x"0023b",
8000=>x"0023b",
8001=>x"0023b",
8002=>x"0023b",
8003=>x"0023b",
8004=>x"0023b",
8005=>x"0023b",
8006=>x"0023b",
8007=>x"0023b",
8008=>x"0023c",
8009=>x"0023c",
8010=>x"0023c",
8011=>x"0023c",
8012=>x"0023c",
8013=>x"0023c",
8014=>x"0023c",
8015=>x"0023c",
8016=>x"0023c",
8017=>x"0023c",
8018=>x"0023c",
8019=>x"0023c",
8020=>x"0023c",
8021=>x"0023c",
8022=>x"0023d",
8023=>x"0023d",
8024=>x"0023d",
8025=>x"0023d",
8026=>x"0023d",
8027=>x"0023d",
8028=>x"0023d",
8029=>x"0023d",
8030=>x"0023d",
8031=>x"0023d",
8032=>x"0023d",
8033=>x"0023d",
8034=>x"0023d",
8035=>x"0023d",
8036=>x"0023e",
8037=>x"0023e",
8038=>x"0023e",
8039=>x"0023e",
8040=>x"0023e",
8041=>x"0023e",
8042=>x"0023e",
8043=>x"0023e",
8044=>x"0023e",
8045=>x"0023e",
8046=>x"0023e",
8047=>x"0023e",
8048=>x"0023e",
8049=>x"0023e",
8050=>x"0023f",
8051=>x"0023f",
8052=>x"0023f",
8053=>x"0023f",
8054=>x"0023f",
8055=>x"0023f",
8056=>x"0023f",
8057=>x"0023f",
8058=>x"0023f",
8059=>x"0023f",
8060=>x"0023f",
8061=>x"0023f",
8062=>x"0023f",
8063=>x"0023f",
8064=>x"00240",
8065=>x"00240",
8066=>x"00240",
8067=>x"00240",
8068=>x"00240",
8069=>x"00240",
8070=>x"00240",
8071=>x"00240",
8072=>x"00240",
8073=>x"00240",
8074=>x"00240",
8075=>x"00240",
8076=>x"00240",
8077=>x"00240",
8078=>x"00241",
8079=>x"00241",
8080=>x"00241",
8081=>x"00241",
8082=>x"00241",
8083=>x"00241",
8084=>x"00241",
8085=>x"00241",
8086=>x"00241",
8087=>x"00241",
8088=>x"00241",
8089=>x"00241",
8090=>x"00241",
8091=>x"00241",
8092=>x"00242",
8093=>x"00242",
8094=>x"00242",
8095=>x"00242",
8096=>x"00242",
8097=>x"00242",
8098=>x"00242",
8099=>x"00242",
8100=>x"00242",
8101=>x"00242",
8102=>x"00242",
8103=>x"00242",
8104=>x"00242",
8105=>x"00242",
8106=>x"00243",
8107=>x"00243",
8108=>x"00243",
8109=>x"00243",
8110=>x"00243",
8111=>x"00243",
8112=>x"00243",
8113=>x"00243",
8114=>x"00243",
8115=>x"00243",
8116=>x"00243",
8117=>x"00243",
8118=>x"00243",
8119=>x"00243",
8120=>x"00244",
8121=>x"00244",
8122=>x"00244",
8123=>x"00244",
8124=>x"00244",
8125=>x"00244",
8126=>x"00244",
8127=>x"00244",
8128=>x"00244",
8129=>x"00244",
8130=>x"00244",
8131=>x"00244",
8132=>x"00244",
8133=>x"00244",
8134=>x"00245",
8135=>x"00245",
8136=>x"00245",
8137=>x"00245",
8138=>x"00245",
8139=>x"00245",
8140=>x"00245",
8141=>x"00245",
8142=>x"00245",
8143=>x"00245",
8144=>x"00245",
8145=>x"00245",
8146=>x"00245",
8147=>x"00245",
8148=>x"00246",
8149=>x"00246",
8150=>x"00246",
8151=>x"00246",
8152=>x"00246",
8153=>x"00246",
8154=>x"00246",
8155=>x"00246",
8156=>x"00246",
8157=>x"00246",
8158=>x"00246",
8159=>x"00246",
8160=>x"00246",
8161=>x"00246",
8162=>x"00247",
8163=>x"00247",
8164=>x"00247",
8165=>x"00247",
8166=>x"00247",
8167=>x"00247",
8168=>x"00247",
8169=>x"00247",
8170=>x"00247",
8171=>x"00247",
8172=>x"00247",
8173=>x"00247",
8174=>x"00247",
8175=>x"00247",
8176=>x"00248",
8177=>x"00248",
8178=>x"00248",
8179=>x"00248",
8180=>x"00248",
8181=>x"00248",
8182=>x"00248",
8183=>x"00248",
8184=>x"00248",
8185=>x"00248",
8186=>x"00248",
8187=>x"00248",
8188=>x"00248",
8189=>x"00248",
8190=>x"00249",
8191=>x"00249",
8192=>x"00249",
8193=>x"00249",
8194=>x"00249",
8195=>x"00249",
8196=>x"00249",
8197=>x"00249",
8198=>x"00249",
8199=>x"00249",
8200=>x"00249",
8201=>x"00249",
8202=>x"00249",
8203=>x"00249",
8204=>x"0024a",
8205=>x"0024a",
8206=>x"0024a",
8207=>x"0024a",
8208=>x"0024a",
8209=>x"0024a",
8210=>x"0024a",
8211=>x"0024a",
8212=>x"0024a",
8213=>x"0024a",
8214=>x"0024a",
8215=>x"0024a",
8216=>x"0024a",
8217=>x"0024a",
8218=>x"0024b",
8219=>x"0024b",
8220=>x"0024b",
8221=>x"0024b",
8222=>x"0024b",
8223=>x"0024b",
8224=>x"0024b",
8225=>x"0024b",
8226=>x"0024b",
8227=>x"0024b",
8228=>x"0024b",
8229=>x"0024b",
8230=>x"0024b",
8231=>x"0024b",
8232=>x"0024c",
8233=>x"0024c",
8234=>x"0024c",
8235=>x"0024c",
8236=>x"0024c",
8237=>x"0024c",
8238=>x"0024c",
8239=>x"0024c",
8240=>x"0024c",
8241=>x"0024c",
8242=>x"0024c",
8243=>x"0024c",
8244=>x"0024c",
8245=>x"0024c",
8246=>x"0024d",
8247=>x"0024d",
8248=>x"0024d",
8249=>x"0024d",
8250=>x"0024d",
8251=>x"0024d",
8252=>x"0024d",
8253=>x"0024d",
8254=>x"0024d",
8255=>x"0024d",
8256=>x"0024d",
8257=>x"0024d",
8258=>x"0024d",
8259=>x"0024d",
8260=>x"0024e",
8261=>x"0024e",
8262=>x"0024e",
8263=>x"0024e",
8264=>x"0024e",
8265=>x"0024e",
8266=>x"0024e",
8267=>x"0024e",
8268=>x"0024e",
8269=>x"0024e",
8270=>x"0024e",
8271=>x"0024e",
8272=>x"0024e",
8273=>x"0024e",
8274=>x"0024f",
8275=>x"0024f",
8276=>x"0024f",
8277=>x"0024f",
8278=>x"0024f",
8279=>x"0024f",
8280=>x"0024f",
8281=>x"0024f",
8282=>x"0024f",
8283=>x"0024f",
8284=>x"0024f",
8285=>x"0024f",
8286=>x"0024f",
8287=>x"0024f",
8288=>x"00250",
8289=>x"00250",
8290=>x"00250",
8291=>x"00250",
8292=>x"00250",
8293=>x"00250",
8294=>x"00250",
8295=>x"00250",
8296=>x"00250",
8297=>x"00250",
8298=>x"00250",
8299=>x"00250",
8300=>x"00250",
8301=>x"00250",
8302=>x"00251",
8303=>x"00251",
8304=>x"00251",
8305=>x"00251",
8306=>x"00251",
8307=>x"00251",
8308=>x"00251",
8309=>x"00251",
8310=>x"00251",
8311=>x"00251",
8312=>x"00251",
8313=>x"00251",
8314=>x"00251",
8315=>x"00251",
8316=>x"00252",
8317=>x"00252",
8318=>x"00252",
8319=>x"00252",
8320=>x"00252",
8321=>x"00252",
8322=>x"00252",
8323=>x"00252",
8324=>x"00252",
8325=>x"00252",
8326=>x"00252",
8327=>x"00252",
8328=>x"00252",
8329=>x"00252",
8330=>x"00253",
8331=>x"00253",
8332=>x"00253",
8333=>x"00253",
8334=>x"00253",
8335=>x"00253",
8336=>x"00253",
8337=>x"00253",
8338=>x"00253",
8339=>x"00253",
8340=>x"00253",
8341=>x"00253",
8342=>x"00253",
8343=>x"00253",
8344=>x"00254",
8345=>x"00254",
8346=>x"00254",
8347=>x"00254",
8348=>x"00254",
8349=>x"00254",
8350=>x"00254",
8351=>x"00254",
8352=>x"00254",
8353=>x"00254",
8354=>x"00254",
8355=>x"00254",
8356=>x"00254",
8357=>x"00254",
8358=>x"00255",
8359=>x"00255",
8360=>x"00255",
8361=>x"00255",
8362=>x"00255",
8363=>x"00255",
8364=>x"00255",
8365=>x"00255",
8366=>x"00255",
8367=>x"00255",
8368=>x"00255",
8369=>x"00255",
8370=>x"00255",
8371=>x"00255",
8372=>x"00256",
8373=>x"00256",
8374=>x"00256",
8375=>x"00256",
8376=>x"00256",
8377=>x"00256",
8378=>x"00256",
8379=>x"00256",
8380=>x"00256",
8381=>x"00256",
8382=>x"00256",
8383=>x"00256",
8384=>x"00256",
8385=>x"00256",
8386=>x"00257",
8387=>x"00257",
8388=>x"00257",
8389=>x"00257",
8390=>x"00257",
8391=>x"00257",
8392=>x"00257",
8393=>x"00257",
8394=>x"00257",
8395=>x"00257",
8396=>x"00257",
8397=>x"00257",
8398=>x"00257",
8399=>x"00257",
8400=>x"00258",
8401=>x"00258",
8402=>x"00258",
8403=>x"00258",
8404=>x"00258",
8405=>x"00258",
8406=>x"00258",
8407=>x"00258",
8408=>x"00258",
8409=>x"00258",
8410=>x"00258",
8411=>x"00258",
8412=>x"00258",
8413=>x"00258",
8414=>x"00259",
8415=>x"00259",
8416=>x"00259",
8417=>x"00259",
8418=>x"00259",
8419=>x"00259",
8420=>x"00259",
8421=>x"00259",
8422=>x"00259",
8423=>x"00259",
8424=>x"00259",
8425=>x"00259",
8426=>x"00259",
8427=>x"00259",
8428=>x"0025a",
8429=>x"0025a",
8430=>x"0025a",
8431=>x"0025a",
8432=>x"0025a",
8433=>x"0025a",
8434=>x"0025a",
8435=>x"0025a",
8436=>x"0025a",
8437=>x"0025a",
8438=>x"0025a",
8439=>x"0025a",
8440=>x"0025a",
8441=>x"0025a",
8442=>x"0025b",
8443=>x"0025b",
8444=>x"0025b",
8445=>x"0025b",
8446=>x"0025b",
8447=>x"0025b",
8448=>x"0025b",
8449=>x"0025b",
8450=>x"0025b",
8451=>x"0025b",
8452=>x"0025b",
8453=>x"0025b",
8454=>x"0025b",
8455=>x"0025b",
8456=>x"0025c",
8457=>x"0025c",
8458=>x"0025c",
8459=>x"0025c",
8460=>x"0025c",
8461=>x"0025c",
8462=>x"0025c",
8463=>x"0025c",
8464=>x"0025c",
8465=>x"0025c",
8466=>x"0025c",
8467=>x"0025c",
8468=>x"0025c",
8469=>x"0025c",
8470=>x"0025d",
8471=>x"0025d",
8472=>x"0025d",
8473=>x"0025d",
8474=>x"0025d",
8475=>x"0025d",
8476=>x"0025d",
8477=>x"0025d",
8478=>x"0025d",
8479=>x"0025d",
8480=>x"0025d",
8481=>x"0025d",
8482=>x"0025d",
8483=>x"0025d",
8484=>x"0025e",
8485=>x"0025e",
8486=>x"0025e",
8487=>x"0025e",
8488=>x"0025e",
8489=>x"0025e",
8490=>x"0025e",
8491=>x"0025e",
8492=>x"0025e",
8493=>x"0025e",
8494=>x"0025e",
8495=>x"0025e",
8496=>x"0025e",
8497=>x"0025e",
8498=>x"0025f",
8499=>x"0025f",
8500=>x"0025f",
8501=>x"0025f",
8502=>x"0025f",
8503=>x"0025f",
8504=>x"0025f",
8505=>x"0025f",
8506=>x"0025f",
8507=>x"0025f",
8508=>x"0025f",
8509=>x"0025f",
8510=>x"0025f",
8511=>x"0025f",
8512=>x"00260",
8513=>x"00260",
8514=>x"00260",
8515=>x"00260",
8516=>x"00260",
8517=>x"00260",
8518=>x"00260",
8519=>x"00260",
8520=>x"00260",
8521=>x"00260",
8522=>x"00260",
8523=>x"00260",
8524=>x"00260",
8525=>x"00260",
8526=>x"00261",
8527=>x"00261",
8528=>x"00261",
8529=>x"00261",
8530=>x"00261",
8531=>x"00261",
8532=>x"00261",
8533=>x"00261",
8534=>x"00261",
8535=>x"00261",
8536=>x"00261",
8537=>x"00261",
8538=>x"00261",
8539=>x"00261",
8540=>x"00262",
8541=>x"00262",
8542=>x"00262",
8543=>x"00262",
8544=>x"00262",
8545=>x"00262",
8546=>x"00262",
8547=>x"00262",
8548=>x"00262",
8549=>x"00262",
8550=>x"00262",
8551=>x"00262",
8552=>x"00262",
8553=>x"00262",
8554=>x"00263",
8555=>x"00263",
8556=>x"00263",
8557=>x"00263",
8558=>x"00263",
8559=>x"00263",
8560=>x"00263",
8561=>x"00263",
8562=>x"00263",
8563=>x"00263",
8564=>x"00263",
8565=>x"00263",
8566=>x"00263",
8567=>x"00263",
8568=>x"00264",
8569=>x"00264",
8570=>x"00264",
8571=>x"00264",
8572=>x"00264",
8573=>x"00264",
8574=>x"00264",
8575=>x"00264",
8576=>x"00264",
8577=>x"00264",
8578=>x"00264",
8579=>x"00264",
8580=>x"00264",
8581=>x"00264",
8582=>x"00265",
8583=>x"00265",
8584=>x"00265",
8585=>x"00265",
8586=>x"00265",
8587=>x"00265",
8588=>x"00265",
8589=>x"00265",
8590=>x"00265",
8591=>x"00265",
8592=>x"00265",
8593=>x"00265",
8594=>x"00265",
8595=>x"00265",
8596=>x"00266",
8597=>x"00266",
8598=>x"00266",
8599=>x"00266",
8600=>x"00266",
8601=>x"00266",
8602=>x"00266",
8603=>x"00266",
8604=>x"00266",
8605=>x"00266",
8606=>x"00266",
8607=>x"00266",
8608=>x"00266",
8609=>x"00266",
8610=>x"00267",
8611=>x"00267",
8612=>x"00267",
8613=>x"00267",
8614=>x"00267",
8615=>x"00267",
8616=>x"00267",
8617=>x"00267",
8618=>x"00267",
8619=>x"00267",
8620=>x"00267",
8621=>x"00267",
8622=>x"00267",
8623=>x"00267",
8624=>x"00268",
8625=>x"00268",
8626=>x"00268",
8627=>x"00268",
8628=>x"00268",
8629=>x"00268",
8630=>x"00268",
8631=>x"00268",
8632=>x"00268",
8633=>x"00268",
8634=>x"00268",
8635=>x"00268",
8636=>x"00268",
8637=>x"00268",
8638=>x"00269",
8639=>x"00269",
8640=>x"00269",
8641=>x"00269",
8642=>x"00269",
8643=>x"00269",
8644=>x"00269",
8645=>x"00269",
8646=>x"00269",
8647=>x"00269",
8648=>x"00269",
8649=>x"00269",
8650=>x"00269",
8651=>x"00269",
8652=>x"0026a",
8653=>x"0026a",
8654=>x"0026a",
8655=>x"0026a",
8656=>x"0026a",
8657=>x"0026a",
8658=>x"0026a",
8659=>x"0026a",
8660=>x"0026a",
8661=>x"0026a",
8662=>x"0026a",
8663=>x"0026a",
8664=>x"0026a",
8665=>x"0026a",
8666=>x"0026b",
8667=>x"0026b",
8668=>x"0026b",
8669=>x"0026b",
8670=>x"0026b",
8671=>x"0026b",
8672=>x"0026b",
8673=>x"0026b",
8674=>x"0026b",
8675=>x"0026b",
8676=>x"0026b",
8677=>x"0026b",
8678=>x"0026b",
8679=>x"0026b",
8680=>x"0026c",
8681=>x"0026c",
8682=>x"0026c",
8683=>x"0026c",
8684=>x"0026c",
8685=>x"0026c",
8686=>x"0026c",
8687=>x"0026c",
8688=>x"0026c",
8689=>x"0026c",
8690=>x"0026c",
8691=>x"0026c",
8692=>x"0026c",
8693=>x"0026c",
8694=>x"0026d",
8695=>x"0026d",
8696=>x"0026d",
8697=>x"0026d",
8698=>x"0026d",
8699=>x"0026d",
8700=>x"0026d",
8701=>x"0026d",
8702=>x"0026d",
8703=>x"0026d",
8704=>x"0026d",
8705=>x"0026d",
8706=>x"0026d",
8707=>x"0026d",
8708=>x"0026e",
8709=>x"0026e",
8710=>x"0026e",
8711=>x"0026e",
8712=>x"0026e",
8713=>x"0026e",
8714=>x"0026e",
8715=>x"0026e",
8716=>x"0026e",
8717=>x"0026e",
8718=>x"0026e",
8719=>x"0026e",
8720=>x"0026e",
8721=>x"0026e",
8722=>x"0026f",
8723=>x"0026f",
8724=>x"0026f",
8725=>x"0026f",
8726=>x"0026f",
8727=>x"0026f",
8728=>x"0026f",
8729=>x"0026f",
8730=>x"0026f",
8731=>x"0026f",
8732=>x"0026f",
8733=>x"0026f",
8734=>x"0026f",
8735=>x"0026f",
8736=>x"00270",
8737=>x"00270",
8738=>x"00270",
8739=>x"00270",
8740=>x"00270",
8741=>x"00270",
8742=>x"00270",
8743=>x"00270",
8744=>x"00270",
8745=>x"00270",
8746=>x"00270",
8747=>x"00270",
8748=>x"00270",
8749=>x"00270",
8750=>x"00271",
8751=>x"00271",
8752=>x"00271",
8753=>x"00271",
8754=>x"00271",
8755=>x"00271",
8756=>x"00271",
8757=>x"00271",
8758=>x"00271",
8759=>x"00271",
8760=>x"00271",
8761=>x"00271",
8762=>x"00271",
8763=>x"00271",
8764=>x"00272",
8765=>x"00272",
8766=>x"00272",
8767=>x"00272",
8768=>x"00272",
8769=>x"00272",
8770=>x"00272",
8771=>x"00272",
8772=>x"00272",
8773=>x"00272",
8774=>x"00272",
8775=>x"00272",
8776=>x"00272",
8777=>x"00272",
8778=>x"00273",
8779=>x"00273",
8780=>x"00273",
8781=>x"00273",
8782=>x"00273",
8783=>x"00273",
8784=>x"00273",
8785=>x"00273",
8786=>x"00273",
8787=>x"00273",
8788=>x"00273",
8789=>x"00273",
8790=>x"00273",
8791=>x"00273",
8792=>x"00274",
8793=>x"00274",
8794=>x"00274",
8795=>x"00274",
8796=>x"00274",
8797=>x"00274",
8798=>x"00274",
8799=>x"00274",
8800=>x"00274",
8801=>x"00274",
8802=>x"00274",
8803=>x"00274",
8804=>x"00274",
8805=>x"00274",
8806=>x"00275",
8807=>x"00275",
8808=>x"00275",
8809=>x"00275",
8810=>x"00275",
8811=>x"00275",
8812=>x"00275",
8813=>x"00275",
8814=>x"00275",
8815=>x"00275",
8816=>x"00275",
8817=>x"00275",
8818=>x"00275",
8819=>x"00275",
8820=>x"00276",
8821=>x"00276",
8822=>x"00276",
8823=>x"00276",
8824=>x"00276",
8825=>x"00276",
8826=>x"00276",
8827=>x"00276",
8828=>x"00276",
8829=>x"00276",
8830=>x"00276",
8831=>x"00276",
8832=>x"00276",
8833=>x"00276",
8834=>x"00277",
8835=>x"00277",
8836=>x"00277",
8837=>x"00277",
8838=>x"00277",
8839=>x"00277",
8840=>x"00277",
8841=>x"00277",
8842=>x"00277",
8843=>x"00277",
8844=>x"00277",
8845=>x"00277",
8846=>x"00277",
8847=>x"00277",
8848=>x"00278",
8849=>x"00278",
8850=>x"00278",
8851=>x"00278",
8852=>x"00278",
8853=>x"00278",
8854=>x"00278",
8855=>x"00278",
8856=>x"00278",
8857=>x"00278",
8858=>x"00278",
8859=>x"00278",
8860=>x"00278",
8861=>x"00278",
8862=>x"00279",
8863=>x"00279",
8864=>x"00279",
8865=>x"00279",
8866=>x"00279",
8867=>x"00279",
8868=>x"00279",
8869=>x"00279",
8870=>x"00279",
8871=>x"00279",
8872=>x"00279",
8873=>x"00279",
8874=>x"00279",
8875=>x"00279",
8876=>x"0027a",
8877=>x"0027a",
8878=>x"0027a",
8879=>x"0027a",
8880=>x"0027a",
8881=>x"0027a",
8882=>x"0027a",
8883=>x"0027a",
8884=>x"0027a",
8885=>x"0027a",
8886=>x"0027a",
8887=>x"0027a",
8888=>x"0027a",
8889=>x"0027a",
8890=>x"0027b",
8891=>x"0027b",
8892=>x"0027b",
8893=>x"0027b",
8894=>x"0027b",
8895=>x"0027b",
8896=>x"0027b",
8897=>x"0027b",
8898=>x"0027b",
8899=>x"0027b",
8900=>x"0027b",
8901=>x"0027b",
8902=>x"0027b",
8903=>x"0027b",
8904=>x"0027c",
8905=>x"0027c",
8906=>x"0027c",
8907=>x"0027c",
8908=>x"0027c",
8909=>x"0027c",
8910=>x"0027c",
8911=>x"0027c",
8912=>x"0027c",
8913=>x"0027c",
8914=>x"0027c",
8915=>x"0027c",
8916=>x"0027c",
8917=>x"0027c",
8918=>x"0027d",
8919=>x"0027d",
8920=>x"0027d",
8921=>x"0027d",
8922=>x"0027d",
8923=>x"0027d",
8924=>x"0027d",
8925=>x"0027d",
8926=>x"0027d",
8927=>x"0027d",
8928=>x"0027d",
8929=>x"0027d",
8930=>x"0027d",
8931=>x"0027d",
8932=>x"0027e",
8933=>x"0027e",
8934=>x"0027e",
8935=>x"0027e",
8936=>x"0027e",
8937=>x"0027e",
8938=>x"0027e",
8939=>x"0027e",
8940=>x"0027e",
8941=>x"0027e",
8942=>x"0027e",
8943=>x"0027e",
8944=>x"0027e",
8945=>x"0027e",
8946=>x"0027f",
8947=>x"0027f",
8948=>x"0027f",
8949=>x"0027f",
8950=>x"0027f",
8951=>x"0027f",
8952=>x"0027f",
8953=>x"0027f",
8954=>x"0027f",
8955=>x"0027f",
8956=>x"0027f",
8957=>x"0027f",
8958=>x"0027f",
8959=>x"0027f",
8960=>x"00280",
8961=>x"00280",
8962=>x"00280",
8963=>x"00280",
8964=>x"00280",
8965=>x"00280",
8966=>x"00280",
8967=>x"00280",
8968=>x"00280",
8969=>x"00280",
8970=>x"00280",
8971=>x"00280",
8972=>x"00280",
8973=>x"00280",
8974=>x"00281",
8975=>x"00281",
8976=>x"00281",
8977=>x"00281",
8978=>x"00281",
8979=>x"00281",
8980=>x"00281",
8981=>x"00281",
8982=>x"00281",
8983=>x"00281",
8984=>x"00281",
8985=>x"00281",
8986=>x"00281",
8987=>x"00281",
8988=>x"00282",
8989=>x"00282",
8990=>x"00282",
8991=>x"00282",
8992=>x"00282",
8993=>x"00282",
8994=>x"00282",
8995=>x"00282",
8996=>x"00282",
8997=>x"00282",
8998=>x"00282",
8999=>x"00282",
9000=>x"00282",
9001=>x"00282",
9002=>x"00283",
9003=>x"00283",
9004=>x"00283",
9005=>x"00283",
9006=>x"00283",
9007=>x"00283",
9008=>x"00283",
9009=>x"00283",
9010=>x"00283",
9011=>x"00283",
9012=>x"00283",
9013=>x"00283",
9014=>x"00283",
9015=>x"00283",
9016=>x"00284",
9017=>x"00284",
9018=>x"00284",
9019=>x"00284",
9020=>x"00284",
9021=>x"00284",
9022=>x"00284",
9023=>x"00284",
9024=>x"00284",
9025=>x"00284",
9026=>x"00284",
9027=>x"00284",
9028=>x"00284",
9029=>x"00284",
9030=>x"00285",
9031=>x"00285",
9032=>x"00285",
9033=>x"00285",
9034=>x"00285",
9035=>x"00285",
9036=>x"00285",
9037=>x"00285",
9038=>x"00285",
9039=>x"00285",
9040=>x"00285",
9041=>x"00285",
9042=>x"00285",
9043=>x"00285",
9044=>x"00286",
9045=>x"00286",
9046=>x"00286",
9047=>x"00286",
9048=>x"00286",
9049=>x"00286",
9050=>x"00286",
9051=>x"00286",
9052=>x"00286",
9053=>x"00286",
9054=>x"00286",
9055=>x"00286",
9056=>x"00286",
9057=>x"00286",
9058=>x"00287",
9059=>x"00287",
9060=>x"00287",
9061=>x"00287",
9062=>x"00287",
9063=>x"00287",
9064=>x"00287",
9065=>x"00287",
9066=>x"00287",
9067=>x"00287",
9068=>x"00287",
9069=>x"00287",
9070=>x"00287",
9071=>x"00287",
9072=>x"00288",
9073=>x"00288",
9074=>x"00288",
9075=>x"00288",
9076=>x"00288",
9077=>x"00288",
9078=>x"00288",
9079=>x"00288",
9080=>x"00288",
9081=>x"00288",
9082=>x"00288",
9083=>x"00288",
9084=>x"00288",
9085=>x"00288",
9086=>x"00289",
9087=>x"00289",
9088=>x"00289",
9089=>x"00289",
9090=>x"00289",
9091=>x"00289",
9092=>x"00289",
9093=>x"00289",
9094=>x"00289",
9095=>x"00289",
9096=>x"00289",
9097=>x"00289",
9098=>x"00289",
9099=>x"00289",
9100=>x"0028a",
9101=>x"0028a",
9102=>x"0028a",
9103=>x"0028a",
9104=>x"0028a",
9105=>x"0028a",
9106=>x"0028a",
9107=>x"0028a",
9108=>x"0028a",
9109=>x"0028a",
9110=>x"0028a",
9111=>x"0028a",
9112=>x"0028a",
9113=>x"0028a",
9114=>x"0028b",
9115=>x"0028b",
9116=>x"0028b",
9117=>x"0028b",
9118=>x"0028b",
9119=>x"0028b",
9120=>x"0028b",
9121=>x"0028b",
9122=>x"0028b",
9123=>x"0028b",
9124=>x"0028b",
9125=>x"0028b",
9126=>x"0028b",
9127=>x"0028b",
9128=>x"0028c",
9129=>x"0028c",
9130=>x"0028c",
9131=>x"0028c",
9132=>x"0028c",
9133=>x"0028c",
9134=>x"0028c",
9135=>x"0028c",
9136=>x"0028c",
9137=>x"0028c",
9138=>x"0028c",
9139=>x"0028c",
9140=>x"0028c",
9141=>x"0028c",
9142=>x"0028d",
9143=>x"0028d",
9144=>x"0028d",
9145=>x"0028d",
9146=>x"0028d",
9147=>x"0028d",
9148=>x"0028d",
9149=>x"0028d",
9150=>x"0028d",
9151=>x"0028d",
9152=>x"0028d",
9153=>x"0028d",
9154=>x"0028d",
9155=>x"0028d",
9156=>x"0028e",
9157=>x"0028e",
9158=>x"0028e",
9159=>x"0028e",
9160=>x"0028e",
9161=>x"0028e",
9162=>x"0028e",
9163=>x"0028e",
9164=>x"0028e",
9165=>x"0028e",
9166=>x"0028e",
9167=>x"0028e",
9168=>x"0028e",
9169=>x"0028e",
9170=>x"0028f",
9171=>x"0028f",
9172=>x"0028f",
9173=>x"0028f",
9174=>x"0028f",
9175=>x"0028f",
9176=>x"0028f",
9177=>x"0028f",
9178=>x"0028f",
9179=>x"0028f",
9180=>x"0028f",
9181=>x"0028f",
9182=>x"0028f",
9183=>x"0028f",
9184=>x"00290",
9185=>x"00290",
9186=>x"00290",
9187=>x"00290",
9188=>x"00290",
9189=>x"00290",
9190=>x"00290",
9191=>x"00290",
9192=>x"00290",
9193=>x"00290",
9194=>x"00290",
9195=>x"00290",
9196=>x"00290",
9197=>x"00290",
9198=>x"00291",
9199=>x"00291",
9200=>x"00291",
9201=>x"00291",
9202=>x"00291",
9203=>x"00291",
9204=>x"00291",
9205=>x"00291",
9206=>x"00291",
9207=>x"00291",
9208=>x"00291",
9209=>x"00291",
9210=>x"00291",
9211=>x"00291",
9212=>x"00292",
9213=>x"00292",
9214=>x"00292",
9215=>x"00292",
9216=>x"00292",
9217=>x"00292",
9218=>x"00292",
9219=>x"00292",
9220=>x"00292",
9221=>x"00292",
9222=>x"00292",
9223=>x"00292",
9224=>x"00292",
9225=>x"00292",
9226=>x"00293",
9227=>x"00293",
9228=>x"00293",
9229=>x"00293",
9230=>x"00293",
9231=>x"00293",
9232=>x"00293",
9233=>x"00293",
9234=>x"00293",
9235=>x"00293",
9236=>x"00293",
9237=>x"00293",
9238=>x"00293",
9239=>x"00293",
9240=>x"00294",
9241=>x"00294",
9242=>x"00294",
9243=>x"00294",
9244=>x"00294",
9245=>x"00294",
9246=>x"00294",
9247=>x"00294",
9248=>x"00294",
9249=>x"00294",
9250=>x"00294",
9251=>x"00294",
9252=>x"00294",
9253=>x"00294",
9254=>x"00295",
9255=>x"00295",
9256=>x"00295",
9257=>x"00295",
9258=>x"00295",
9259=>x"00295",
9260=>x"00295",
9261=>x"00295",
9262=>x"00295",
9263=>x"00295",
9264=>x"00295",
9265=>x"00295",
9266=>x"00295",
9267=>x"00295",
9268=>x"00296",
9269=>x"00296",
9270=>x"00296",
9271=>x"00296",
9272=>x"00296",
9273=>x"00296",
9274=>x"00296",
9275=>x"00296",
9276=>x"00296",
9277=>x"00296",
9278=>x"00296",
9279=>x"00296",
9280=>x"00296",
9281=>x"00296",
9282=>x"00297",
9283=>x"00297",
9284=>x"00297",
9285=>x"00297",
9286=>x"00297",
9287=>x"00297",
9288=>x"00297",
9289=>x"00297",
9290=>x"00297",
9291=>x"00297",
9292=>x"00297",
9293=>x"00297",
9294=>x"00297",
9295=>x"00297",
9296=>x"00298",
9297=>x"00298",
9298=>x"00298",
9299=>x"00298",
9300=>x"00298",
9301=>x"00298",
9302=>x"00298",
9303=>x"00298",
9304=>x"00298",
9305=>x"00298",
9306=>x"00298",
9307=>x"00298",
9308=>x"00298",
9309=>x"00298",
9310=>x"00299",
9311=>x"00299",
9312=>x"00299",
9313=>x"00299",
9314=>x"00299",
9315=>x"00299",
9316=>x"00299",
9317=>x"00299",
9318=>x"00299",
9319=>x"00299",
9320=>x"00299",
9321=>x"00299",
9322=>x"00299",
9323=>x"00299",
9324=>x"0029a",
9325=>x"0029a",
9326=>x"0029a",
9327=>x"0029a",
9328=>x"0029a",
9329=>x"0029a",
9330=>x"0029a",
9331=>x"0029a",
9332=>x"0029a",
9333=>x"0029a",
9334=>x"0029a",
9335=>x"0029a",
9336=>x"0029a",
9337=>x"0029a",
9338=>x"0029b",
9339=>x"0029b",
9340=>x"0029b",
9341=>x"0029b",
9342=>x"0029b",
9343=>x"0029b",
9344=>x"0029b",
9345=>x"0029b",
9346=>x"0029b",
9347=>x"0029b",
9348=>x"0029b",
9349=>x"0029b",
9350=>x"0029b",
9351=>x"0029b",
9352=>x"0029c",
9353=>x"0029c",
9354=>x"0029c",
9355=>x"0029c",
9356=>x"0029c",
9357=>x"0029c",
9358=>x"0029c",
9359=>x"0029c",
9360=>x"0029c",
9361=>x"0029c",
9362=>x"0029c",
9363=>x"0029c",
9364=>x"0029c",
9365=>x"0029c",
9366=>x"0029d",
9367=>x"0029d",
9368=>x"0029d",
9369=>x"0029d",
9370=>x"0029d",
9371=>x"0029d",
9372=>x"0029d",
9373=>x"0029d",
9374=>x"0029d",
9375=>x"0029d",
9376=>x"0029d",
9377=>x"0029d",
9378=>x"0029d",
9379=>x"0029d",
9380=>x"0029e",
9381=>x"0029e",
9382=>x"0029e",
9383=>x"0029e",
9384=>x"0029e",
9385=>x"0029e",
9386=>x"0029e",
9387=>x"0029e",
9388=>x"0029e",
9389=>x"0029e",
9390=>x"0029e",
9391=>x"0029e",
9392=>x"0029e",
9393=>x"0029e",
9394=>x"0029f",
9395=>x"0029f",
9396=>x"0029f",
9397=>x"0029f",
9398=>x"0029f",
9399=>x"0029f",
9400=>x"0029f",
9401=>x"0029f",
9402=>x"0029f",
9403=>x"0029f",
9404=>x"0029f",
9405=>x"0029f",
9406=>x"0029f",
9407=>x"0029f",
9408=>x"002a0",
9409=>x"002a0",
9410=>x"002a0",
9411=>x"002a0",
9412=>x"002a0",
9413=>x"002a0",
9414=>x"002a0",
9415=>x"002a0",
9416=>x"002a0",
9417=>x"002a0",
9418=>x"002a0",
9419=>x"002a0",
9420=>x"002a0",
9421=>x"002a0",
9422=>x"002a1",
9423=>x"002a1",
9424=>x"002a1",
9425=>x"002a1",
9426=>x"002a1",
9427=>x"002a1",
9428=>x"002a1",
9429=>x"002a1",
9430=>x"002a1",
9431=>x"002a1",
9432=>x"002a1",
9433=>x"002a1",
9434=>x"002a1",
9435=>x"002a1",
9436=>x"002a2",
9437=>x"002a2",
9438=>x"002a2",
9439=>x"002a2",
9440=>x"002a2",
9441=>x"002a2",
9442=>x"002a2",
9443=>x"002a2",
9444=>x"002a2",
9445=>x"002a2",
9446=>x"002a2",
9447=>x"002a2",
9448=>x"002a2",
9449=>x"002a2",
9450=>x"002a3",
9451=>x"002a3",
9452=>x"002a3",
9453=>x"002a3",
9454=>x"002a3",
9455=>x"002a3",
9456=>x"002a3",
9457=>x"002a3",
9458=>x"002a3",
9459=>x"002a3",
9460=>x"002a3",
9461=>x"002a3",
9462=>x"002a3",
9463=>x"002a3",
9464=>x"002a4",
9465=>x"002a4",
9466=>x"002a4",
9467=>x"002a4",
9468=>x"002a4",
9469=>x"002a4",
9470=>x"002a4",
9471=>x"002a4",
9472=>x"002a4",
9473=>x"002a4",
9474=>x"002a4",
9475=>x"002a4",
9476=>x"002a4",
9477=>x"002a4",
9478=>x"002a5",
9479=>x"002a5",
9480=>x"002a5",
9481=>x"002a5",
9482=>x"002a5",
9483=>x"002a5",
9484=>x"002a5",
9485=>x"002a5",
9486=>x"002a5",
9487=>x"002a5",
9488=>x"002a5",
9489=>x"002a5",
9490=>x"002a5",
9491=>x"002a5",
9492=>x"002a6",
9493=>x"002a6",
9494=>x"002a6",
9495=>x"002a6",
9496=>x"002a6",
9497=>x"002a6",
9498=>x"002a6",
9499=>x"002a6",
9500=>x"002a6",
9501=>x"002a6",
9502=>x"002a6",
9503=>x"002a6",
9504=>x"002a6",
9505=>x"002a6",
9506=>x"002a7",
9507=>x"002a7",
9508=>x"002a7",
9509=>x"002a7",
9510=>x"002a7",
9511=>x"002a7",
9512=>x"002a7",
9513=>x"002a7",
9514=>x"002a7",
9515=>x"002a7",
9516=>x"002a7",
9517=>x"002a7",
9518=>x"002a7",
9519=>x"002a7",
9520=>x"002a8",
9521=>x"002a8",
9522=>x"002a8",
9523=>x"002a8",
9524=>x"002a8",
9525=>x"002a8",
9526=>x"002a8",
9527=>x"002a8",
9528=>x"002a8",
9529=>x"002a8",
9530=>x"002a8",
9531=>x"002a8",
9532=>x"002a8",
9533=>x"002a8",
9534=>x"002a9",
9535=>x"002a9",
9536=>x"002a9",
9537=>x"002a9",
9538=>x"002a9",
9539=>x"002a9",
9540=>x"002a9",
9541=>x"002a9",
9542=>x"002a9",
9543=>x"002a9",
9544=>x"002a9",
9545=>x"002a9",
9546=>x"002a9",
9547=>x"002a9",
9548=>x"002aa",
9549=>x"002aa",
9550=>x"002aa",
9551=>x"002aa",
9552=>x"002aa",
9553=>x"002aa",
9554=>x"002aa",
9555=>x"002aa",
9556=>x"002aa",
9557=>x"002aa",
9558=>x"002aa",
9559=>x"002aa",
9560=>x"002aa",
9561=>x"002aa",
9562=>x"002ab",
9563=>x"002ab",
9564=>x"002ab",
9565=>x"002ab",
9566=>x"002ab",
9567=>x"002ab",
9568=>x"002ab",
9569=>x"002ab",
9570=>x"002ab",
9571=>x"002ab",
9572=>x"002ab",
9573=>x"002ab",
9574=>x"002ab",
9575=>x"002ab",
9576=>x"002ac",
9577=>x"002ac",
9578=>x"002ac",
9579=>x"002ac",
9580=>x"002ac",
9581=>x"002ac",
9582=>x"002ac",
9583=>x"002ac",
9584=>x"002ac",
9585=>x"002ac",
9586=>x"002ac",
9587=>x"002ac",
9588=>x"002ac",
9589=>x"002ac",
9590=>x"002ad",
9591=>x"002ad",
9592=>x"002ad",
9593=>x"002ad",
9594=>x"002ad",
9595=>x"002ad",
9596=>x"002ad",
9597=>x"002ad",
9598=>x"002ad",
9599=>x"002ad",
9600=>x"002ad",
9601=>x"002ad",
9602=>x"002ad",
9603=>x"002ad",
9604=>x"002ae",
9605=>x"002ae",
9606=>x"002ae",
9607=>x"002ae",
9608=>x"002ae",
9609=>x"002ae",
9610=>x"002ae",
9611=>x"002ae",
9612=>x"002ae",
9613=>x"002ae",
9614=>x"002ae",
9615=>x"002ae",
9616=>x"002ae",
9617=>x"002ae",
9618=>x"002af",
9619=>x"002af",
9620=>x"002af",
9621=>x"002af",
9622=>x"002af",
9623=>x"002af",
9624=>x"002af",
9625=>x"002af",
9626=>x"002af",
9627=>x"002af",
9628=>x"002af",
9629=>x"002af",
9630=>x"002af",
9631=>x"002af",
9632=>x"002b0",
9633=>x"002b0",
9634=>x"002b0",
9635=>x"002b0",
9636=>x"002b0",
9637=>x"002b0",
9638=>x"002b0",
9639=>x"002b0",
9640=>x"002b0",
9641=>x"002b0",
9642=>x"002b0",
9643=>x"002b0",
9644=>x"002b0",
9645=>x"002b0",
9646=>x"002b1",
9647=>x"002b1",
9648=>x"002b1",
9649=>x"002b1",
9650=>x"002b1",
9651=>x"002b1",
9652=>x"002b1",
9653=>x"002b1",
9654=>x"002b1",
9655=>x"002b1",
9656=>x"002b1",
9657=>x"002b1",
9658=>x"002b1",
9659=>x"002b1",
9660=>x"002b2",
9661=>x"002b2",
9662=>x"002b2",
9663=>x"002b2",
9664=>x"002b2",
9665=>x"002b2",
9666=>x"002b2",
9667=>x"002b2",
9668=>x"002b2",
9669=>x"002b2",
9670=>x"002b2",
9671=>x"002b2",
9672=>x"002b2",
9673=>x"002b2",
9674=>x"002b3",
9675=>x"002b3",
9676=>x"002b3",
9677=>x"002b3",
9678=>x"002b3",
9679=>x"002b3",
9680=>x"002b3",
9681=>x"002b3",
9682=>x"002b3",
9683=>x"002b3",
9684=>x"002b3",
9685=>x"002b3",
9686=>x"002b3",
9687=>x"002b3",
9688=>x"002b4",
9689=>x"002b4",
9690=>x"002b4",
9691=>x"002b4",
9692=>x"002b4",
9693=>x"002b4",
9694=>x"002b4",
9695=>x"002b4",
9696=>x"002b4",
9697=>x"002b4",
9698=>x"002b4",
9699=>x"002b4",
9700=>x"002b4",
9701=>x"002b4",
9702=>x"002b5",
9703=>x"002b5",
9704=>x"002b5",
9705=>x"002b5",
9706=>x"002b5",
9707=>x"002b5",
9708=>x"002b5",
9709=>x"002b5",
9710=>x"002b5",
9711=>x"002b5",
9712=>x"002b5",
9713=>x"002b5",
9714=>x"002b5",
9715=>x"002b5",
9716=>x"002b6",
9717=>x"002b6",
9718=>x"002b6",
9719=>x"002b6",
9720=>x"002b6",
9721=>x"002b6",
9722=>x"002b6",
9723=>x"002b6",
9724=>x"002b6",
9725=>x"002b6",
9726=>x"002b6",
9727=>x"002b6",
9728=>x"002b6",
9729=>x"002b6",
9730=>x"002b7",
9731=>x"002b7",
9732=>x"002b7",
9733=>x"002b7",
9734=>x"002b7",
9735=>x"002b7",
9736=>x"002b7",
9737=>x"002b7",
9738=>x"002b7",
9739=>x"002b7",
9740=>x"002b7",
9741=>x"002b7",
9742=>x"002b7",
9743=>x"002b7",
9744=>x"002b8",
9745=>x"002b8",
9746=>x"002b8",
9747=>x"002b8",
9748=>x"002b8",
9749=>x"002b8",
9750=>x"002b8",
9751=>x"002b8",
9752=>x"002b8",
9753=>x"002b8",
9754=>x"002b8",
9755=>x"002b8",
9756=>x"002b8",
9757=>x"002b8",
9758=>x"002b9",
9759=>x"002b9",
9760=>x"002b9",
9761=>x"002b9",
9762=>x"002b9",
9763=>x"002b9",
9764=>x"002b9",
9765=>x"002b9",
9766=>x"002b9",
9767=>x"002b9",
9768=>x"002b9",
9769=>x"002b9",
9770=>x"002b9",
9771=>x"002b9",
9772=>x"002ba",
9773=>x"002ba",
9774=>x"002ba",
9775=>x"002ba",
9776=>x"002ba",
9777=>x"002ba",
9778=>x"002ba",
9779=>x"002ba",
9780=>x"002ba",
9781=>x"002ba",
9782=>x"002ba",
9783=>x"002ba",
9784=>x"002ba",
9785=>x"002ba",
9786=>x"002bb",
9787=>x"002bb",
9788=>x"002bb",
9789=>x"002bb",
9790=>x"002bb",
9791=>x"002bb",
9792=>x"002bb",
9793=>x"002bb",
9794=>x"002bb",
9795=>x"002bb",
9796=>x"002bb",
9797=>x"002bb",
9798=>x"002bb",
9799=>x"002bb",
9800=>x"002bc",
9801=>x"002bc",
9802=>x"002bc",
9803=>x"002bc",
9804=>x"002bc",
9805=>x"002bc",
9806=>x"002bc",
9807=>x"002bc",
9808=>x"002bc",
9809=>x"002bc",
9810=>x"002bc",
9811=>x"002bc",
9812=>x"002bc",
9813=>x"002bc",
9814=>x"002bd",
9815=>x"002bd",
9816=>x"002bd",
9817=>x"002bd",
9818=>x"002bd",
9819=>x"002bd",
9820=>x"002bd",
9821=>x"002bd",
9822=>x"002bd",
9823=>x"002bd",
9824=>x"002bd",
9825=>x"002bd",
9826=>x"002bd",
9827=>x"002bd",
9828=>x"002be",
9829=>x"002be",
9830=>x"002be",
9831=>x"002be",
9832=>x"002be",
9833=>x"002be",
9834=>x"002be",
9835=>x"002be",
9836=>x"002be",
9837=>x"002be",
9838=>x"002be",
9839=>x"002be",
9840=>x"002be",
9841=>x"002be",
9842=>x"002bf",
9843=>x"002bf",
9844=>x"002bf",
9845=>x"002bf",
9846=>x"002bf",
9847=>x"002bf",
9848=>x"002bf",
9849=>x"002bf",
9850=>x"002bf",
9851=>x"002bf",
9852=>x"002bf",
9853=>x"002bf",
9854=>x"002bf",
9855=>x"002bf",
9856=>x"002c0",
9857=>x"002c0",
9858=>x"002c0",
9859=>x"002c0",
9860=>x"002c0",
9861=>x"002c0",
9862=>x"002c0",
9863=>x"002c0",
9864=>x"002c0",
9865=>x"002c0",
9866=>x"002c0",
9867=>x"002c0",
9868=>x"002c0",
9869=>x"002c0",
9870=>x"002c1",
9871=>x"002c1",
9872=>x"002c1",
9873=>x"002c1",
9874=>x"002c1",
9875=>x"002c1",
9876=>x"002c1",
9877=>x"002c1",
9878=>x"002c1",
9879=>x"002c1",
9880=>x"002c1",
9881=>x"002c1",
9882=>x"002c1",
9883=>x"002c1",
9884=>x"002c2",
9885=>x"002c2",
9886=>x"002c2",
9887=>x"002c2",
9888=>x"002c2",
9889=>x"002c2",
9890=>x"002c2",
9891=>x"002c2",
9892=>x"002c2",
9893=>x"002c2",
9894=>x"002c2",
9895=>x"002c2",
9896=>x"002c2",
9897=>x"002c2",
9898=>x"002c3",
9899=>x"002c3",
9900=>x"002c3",
9901=>x"002c3",
9902=>x"002c3",
9903=>x"002c3",
9904=>x"002c3",
9905=>x"002c3",
9906=>x"002c3",
9907=>x"002c3",
9908=>x"002c3",
9909=>x"002c3",
9910=>x"002c3",
9911=>x"002c3",
9912=>x"002c4",
9913=>x"002c4",
9914=>x"002c4",
9915=>x"002c4",
9916=>x"002c4",
9917=>x"002c4",
9918=>x"002c4",
9919=>x"002c4",
9920=>x"002c4",
9921=>x"002c4",
9922=>x"002c4",
9923=>x"002c4",
9924=>x"002c4",
9925=>x"002c4",
9926=>x"002c5",
9927=>x"002c5",
9928=>x"002c5",
9929=>x"002c5",
9930=>x"002c5",
9931=>x"002c5",
9932=>x"002c5",
9933=>x"002c5",
9934=>x"002c5",
9935=>x"002c5",
9936=>x"002c5",
9937=>x"002c5",
9938=>x"002c5",
9939=>x"002c5",
9940=>x"002c6",
9941=>x"002c6",
9942=>x"002c6",
9943=>x"002c6",
9944=>x"002c6",
9945=>x"002c6",
9946=>x"002c6",
9947=>x"002c6",
9948=>x"002c6",
9949=>x"002c6",
9950=>x"002c6",
9951=>x"002c6",
9952=>x"002c6",
9953=>x"002c6",
9954=>x"002c7",
9955=>x"002c7",
9956=>x"002c7",
9957=>x"002c7",
9958=>x"002c7",
9959=>x"002c7",
9960=>x"002c7",
9961=>x"002c7",
9962=>x"002c7",
9963=>x"002c7",
9964=>x"002c7",
9965=>x"002c7",
9966=>x"002c7",
9967=>x"002c7",
9968=>x"002c8",
9969=>x"002c8",
9970=>x"002c8",
9971=>x"002c8",
9972=>x"002c8",
9973=>x"002c8",
9974=>x"002c8",
9975=>x"002c8",
9976=>x"002c8",
9977=>x"002c8",
9978=>x"002c8",
9979=>x"002c8",
9980=>x"002c8",
9981=>x"002c8",
9982=>x"002c9",
9983=>x"002c9",
9984=>x"002c9",
9985=>x"002c9",
9986=>x"002c9",
9987=>x"002c9",
9988=>x"002c9",
9989=>x"002c9",
9990=>x"002c9",
9991=>x"002c9",
9992=>x"002c9",
9993=>x"002c9",
9994=>x"002c9",
9995=>x"002c9",
9996=>x"002ca",
9997=>x"002ca",
9998=>x"002ca",
9999=>x"002ca",
10000=>x"002ca",
10001=>x"002ca",
10002=>x"002ca",
10003=>x"002ca",
10004=>x"002ca",
10005=>x"002ca",
10006=>x"002ca",
10007=>x"002ca",
10008=>x"002ca",
10009=>x"002ca",
10010=>x"002cb",
10011=>x"002cb",
10012=>x"002cb",
10013=>x"002cb",
10014=>x"002cb",
10015=>x"002cb",
10016=>x"002cb",
10017=>x"002cb",
10018=>x"002cb",
10019=>x"002cb",
10020=>x"002cb",
10021=>x"002cb",
10022=>x"002cb",
10023=>x"002cb",
10024=>x"002cc",
10025=>x"002cc",
10026=>x"002cc",
10027=>x"002cc",
10028=>x"002cc",
10029=>x"002cc",
10030=>x"002cc",
10031=>x"002cc",
10032=>x"002cc",
10033=>x"002cc",
10034=>x"002cc",
10035=>x"002cc",
10036=>x"002cc",
10037=>x"002cc",
10038=>x"002cd",
10039=>x"002cd",
10040=>x"002cd",
10041=>x"002cd",
10042=>x"002cd",
10043=>x"002cd",
10044=>x"002cd",
10045=>x"002cd",
10046=>x"002cd",
10047=>x"002cd",
10048=>x"002cd",
10049=>x"002cd",
10050=>x"002cd",
10051=>x"002cd",
10052=>x"002ce",
10053=>x"002ce",
10054=>x"002ce",
10055=>x"002ce",
10056=>x"002ce",
10057=>x"002ce",
10058=>x"002ce",
10059=>x"002ce",
10060=>x"002ce",
10061=>x"002ce",
10062=>x"002ce",
10063=>x"002ce",
10064=>x"002ce",
10065=>x"002ce",
10066=>x"002cf",
10067=>x"002cf",
10068=>x"002cf",
10069=>x"002cf",
10070=>x"002cf",
10071=>x"002cf",
10072=>x"002cf",
10073=>x"002cf",
10074=>x"002cf",
10075=>x"002cf",
10076=>x"002cf",
10077=>x"002cf",
10078=>x"002cf",
10079=>x"002cf",
10080=>x"002d0",
10081=>x"002d0",
10082=>x"002d0",
10083=>x"002d0",
10084=>x"002d0",
10085=>x"002d0",
10086=>x"002d0",
10087=>x"002d0",
10088=>x"002d0",
10089=>x"002d0",
10090=>x"002d0",
10091=>x"002d0",
10092=>x"002d0",
10093=>x"002d0",
10094=>x"002d1",
10095=>x"002d1",
10096=>x"002d1",
10097=>x"002d1",
10098=>x"002d1",
10099=>x"002d1",
10100=>x"002d1",
10101=>x"002d1",
10102=>x"002d1",
10103=>x"002d1",
10104=>x"002d1",
10105=>x"002d1",
10106=>x"002d1",
10107=>x"002d1",
10108=>x"002d2",
10109=>x"002d2",
10110=>x"002d2",
10111=>x"002d2",
10112=>x"002d2",
10113=>x"002d2",
10114=>x"002d2",
10115=>x"002d2",
10116=>x"002d2",
10117=>x"002d2",
10118=>x"002d2",
10119=>x"002d2",
10120=>x"002d2",
10121=>x"002d2",
10122=>x"002d3",
10123=>x"002d3",
10124=>x"002d3",
10125=>x"002d3",
10126=>x"002d3",
10127=>x"002d3",
10128=>x"002d3",
10129=>x"002d3",
10130=>x"002d3",
10131=>x"002d3",
10132=>x"002d3",
10133=>x"002d3",
10134=>x"002d3",
10135=>x"002d3",
10136=>x"002d4",
10137=>x"002d4",
10138=>x"002d4",
10139=>x"002d4",
10140=>x"002d4",
10141=>x"002d4",
10142=>x"002d4",
10143=>x"002d4",
10144=>x"002d4",
10145=>x"002d4",
10146=>x"002d4",
10147=>x"002d4",
10148=>x"002d4",
10149=>x"002d4",
10150=>x"002d5",
10151=>x"002d5",
10152=>x"002d5",
10153=>x"002d5",
10154=>x"002d5",
10155=>x"002d5",
10156=>x"002d5",
10157=>x"002d5",
10158=>x"002d5",
10159=>x"002d5",
10160=>x"002d5",
10161=>x"002d5",
10162=>x"002d5",
10163=>x"002d5",
10164=>x"002d6",
10165=>x"002d6",
10166=>x"002d6",
10167=>x"002d6",
10168=>x"002d6",
10169=>x"002d6",
10170=>x"002d6",
10171=>x"002d6",
10172=>x"002d6",
10173=>x"002d6",
10174=>x"002d6",
10175=>x"002d6",
10176=>x"002d6",
10177=>x"002d6",
10178=>x"002d7",
10179=>x"002d7",
10180=>x"002d7",
10181=>x"002d7",
10182=>x"002d7",
10183=>x"002d7",
10184=>x"002d7",
10185=>x"002d7",
10186=>x"002d7",
10187=>x"002d7",
10188=>x"002d7",
10189=>x"002d7",
10190=>x"002d7",
10191=>x"002d7",
10192=>x"002d8",
10193=>x"002d8",
10194=>x"002d8",
10195=>x"002d8",
10196=>x"002d8",
10197=>x"002d8",
10198=>x"002d8",
10199=>x"002d8",
10200=>x"002d8",
10201=>x"002d8",
10202=>x"002d8",
10203=>x"002d8",
10204=>x"002d8",
10205=>x"002d8",
10206=>x"002d9",
10207=>x"002d9",
10208=>x"002d9",
10209=>x"002d9",
10210=>x"002d9",
10211=>x"002d9",
10212=>x"002d9",
10213=>x"002d9",
10214=>x"002d9",
10215=>x"002d9",
10216=>x"002d9",
10217=>x"002d9",
10218=>x"002d9",
10219=>x"002d9",
10220=>x"002da",
10221=>x"002da",
10222=>x"002da",
10223=>x"002da",
10224=>x"002da",
10225=>x"002da",
10226=>x"002da",
10227=>x"002da",
10228=>x"002da",
10229=>x"002da",
10230=>x"002da",
10231=>x"002da",
10232=>x"002da",
10233=>x"002da",
10234=>x"002db",
10235=>x"002db",
10236=>x"002db",
10237=>x"002db",
10238=>x"002db",
10239=>x"002db",
10240=>x"002db",
10241=>x"002db",
10242=>x"002db",
10243=>x"002db",
10244=>x"002db",
10245=>x"002db",
10246=>x"002db",
10247=>x"002db",
10248=>x"002dc",
10249=>x"002dc",
10250=>x"002dc",
10251=>x"002dc",
10252=>x"002dc",
10253=>x"002dc",
10254=>x"002dc",
10255=>x"002dc",
10256=>x"002dc",
10257=>x"002dc",
10258=>x"002dc",
10259=>x"002dc",
10260=>x"002dc",
10261=>x"002dc",
10262=>x"002dd",
10263=>x"002dd",
10264=>x"002dd",
10265=>x"002dd",
10266=>x"002dd",
10267=>x"002dd",
10268=>x"002dd",
10269=>x"002dd",
10270=>x"002dd",
10271=>x"002dd",
10272=>x"002dd",
10273=>x"002dd",
10274=>x"002dd",
10275=>x"002dd",
10276=>x"002de",
10277=>x"002de",
10278=>x"002de",
10279=>x"002de",
10280=>x"002de",
10281=>x"002de",
10282=>x"002de",
10283=>x"002de",
10284=>x"002de",
10285=>x"002de",
10286=>x"002de",
10287=>x"002de",
10288=>x"002de",
10289=>x"002de",
10290=>x"002df",
10291=>x"002df",
10292=>x"002df",
10293=>x"002df",
10294=>x"002df",
10295=>x"002df",
10296=>x"002df",
10297=>x"002df",
10298=>x"002df",
10299=>x"002df",
10300=>x"002df",
10301=>x"002df",
10302=>x"002df",
10303=>x"002df",
10304=>x"002e0",
10305=>x"002e0",
10306=>x"002e0",
10307=>x"002e0",
10308=>x"002e0",
10309=>x"002e0",
10310=>x"002e0",
10311=>x"002e0",
10312=>x"002e0",
10313=>x"002e0",
10314=>x"002e0",
10315=>x"002e0",
10316=>x"002e0",
10317=>x"002e0",
10318=>x"002e1",
10319=>x"002e1",
10320=>x"002e1",
10321=>x"002e1",
10322=>x"002e1",
10323=>x"002e1",
10324=>x"002e1",
10325=>x"002e1",
10326=>x"002e1",
10327=>x"002e1",
10328=>x"002e1",
10329=>x"002e1",
10330=>x"002e1",
10331=>x"002e1",
10332=>x"002e2",
10333=>x"002e2",
10334=>x"002e2",
10335=>x"002e2",
10336=>x"002e2",
10337=>x"002e2",
10338=>x"002e2",
10339=>x"002e2",
10340=>x"002e2",
10341=>x"002e2",
10342=>x"002e2",
10343=>x"002e2",
10344=>x"002e2",
10345=>x"002e2",
10346=>x"002e3",
10347=>x"002e3",
10348=>x"002e3",
10349=>x"002e3",
10350=>x"002e3",
10351=>x"002e3",
10352=>x"002e3",
10353=>x"002e3",
10354=>x"002e3",
10355=>x"002e3",
10356=>x"002e3",
10357=>x"002e3",
10358=>x"002e3",
10359=>x"002e3",
10360=>x"002e4",
10361=>x"002e4",
10362=>x"002e4",
10363=>x"002e4",
10364=>x"002e4",
10365=>x"002e4",
10366=>x"002e4",
10367=>x"002e4",
10368=>x"002e4",
10369=>x"002e4",
10370=>x"002e4",
10371=>x"002e4",
10372=>x"002e4",
10373=>x"002e4",
10374=>x"002e5",
10375=>x"002e5",
10376=>x"002e5",
10377=>x"002e5",
10378=>x"002e5",
10379=>x"002e5",
10380=>x"002e5",
10381=>x"002e5",
10382=>x"002e5",
10383=>x"002e5",
10384=>x"002e5",
10385=>x"002e5",
10386=>x"002e5",
10387=>x"002e5",
10388=>x"002e6",
10389=>x"002e6",
10390=>x"002e6",
10391=>x"002e6",
10392=>x"002e6",
10393=>x"002e6",
10394=>x"002e6",
10395=>x"002e6",
10396=>x"002e6",
10397=>x"002e6",
10398=>x"002e6",
10399=>x"002e6",
10400=>x"002e6",
10401=>x"002e6",
10402=>x"002e7",
10403=>x"002e7",
10404=>x"002e7",
10405=>x"002e7",
10406=>x"002e7",
10407=>x"002e7",
10408=>x"002e7",
10409=>x"002e7",
10410=>x"002e7",
10411=>x"002e7",
10412=>x"002e7",
10413=>x"002e7",
10414=>x"002e7",
10415=>x"002e7",
10416=>x"002e8",
10417=>x"002e8",
10418=>x"002e8",
10419=>x"002e8",
10420=>x"002e8",
10421=>x"002e8",
10422=>x"002e8",
10423=>x"002e8",
10424=>x"002e8",
10425=>x"002e8",
10426=>x"002e8",
10427=>x"002e8",
10428=>x"002e8",
10429=>x"002e8",
10430=>x"002e9",
10431=>x"002e9",
10432=>x"002e9",
10433=>x"002e9",
10434=>x"002e9",
10435=>x"002e9",
10436=>x"002e9",
10437=>x"002e9",
10438=>x"002e9",
10439=>x"002e9",
10440=>x"002e9",
10441=>x"002e9",
10442=>x"002e9",
10443=>x"002e9",
10444=>x"002ea",
10445=>x"002ea",
10446=>x"002ea",
10447=>x"002ea",
10448=>x"002ea",
10449=>x"002ea",
10450=>x"002ea",
10451=>x"002ea",
10452=>x"002ea",
10453=>x"002ea",
10454=>x"002ea",
10455=>x"002ea",
10456=>x"002ea",
10457=>x"002ea",
10458=>x"002eb",
10459=>x"002eb",
10460=>x"002eb",
10461=>x"002eb",
10462=>x"002eb",
10463=>x"002eb",
10464=>x"002eb",
10465=>x"002eb",
10466=>x"002eb",
10467=>x"002eb",
10468=>x"002eb",
10469=>x"002eb",
10470=>x"002eb",
10471=>x"002eb",
10472=>x"002ec",
10473=>x"002ec",
10474=>x"002ec",
10475=>x"002ec",
10476=>x"002ec",
10477=>x"002ec",
10478=>x"002ec",
10479=>x"002ec",
10480=>x"002ec",
10481=>x"002ec",
10482=>x"002ec",
10483=>x"002ec",
10484=>x"002ec",
10485=>x"002ec",
10486=>x"002ed",
10487=>x"002ed",
10488=>x"002ed",
10489=>x"002ed",
10490=>x"002ed",
10491=>x"002ed",
10492=>x"002ed",
10493=>x"002ed",
10494=>x"002ed",
10495=>x"002ed",
10496=>x"002ed",
10497=>x"002ed",
10498=>x"002ed",
10499=>x"002ed",
10500=>x"002ee",
10501=>x"002ee",
10502=>x"002ee",
10503=>x"002ee",
10504=>x"002ee",
10505=>x"002ee",
10506=>x"002ee",
10507=>x"002ee",
10508=>x"002ee",
10509=>x"002ee",
10510=>x"002ee",
10511=>x"002ee",
10512=>x"002ee",
10513=>x"002ee",
10514=>x"002ef",
10515=>x"002ef",
10516=>x"002ef",
10517=>x"002ef",
10518=>x"002ef",
10519=>x"002ef",
10520=>x"002ef",
10521=>x"002ef",
10522=>x"002ef",
10523=>x"002ef",
10524=>x"002ef",
10525=>x"002ef",
10526=>x"002ef",
10527=>x"002ef",
10528=>x"002f0",
10529=>x"002f0",
10530=>x"002f0",
10531=>x"002f0",
10532=>x"002f0",
10533=>x"002f0",
10534=>x"002f0",
10535=>x"002f0",
10536=>x"002f0",
10537=>x"002f0",
10538=>x"002f0",
10539=>x"002f0",
10540=>x"002f0",
10541=>x"002f0",
10542=>x"002f1",
10543=>x"002f1",
10544=>x"002f1",
10545=>x"002f1",
10546=>x"002f1",
10547=>x"002f1",
10548=>x"002f1",
10549=>x"002f1",
10550=>x"002f1",
10551=>x"002f1",
10552=>x"002f1",
10553=>x"002f1",
10554=>x"002f1",
10555=>x"002f1",
10556=>x"002f2",
10557=>x"002f2",
10558=>x"002f2",
10559=>x"002f2",
10560=>x"002f2",
10561=>x"002f2",
10562=>x"002f2",
10563=>x"002f2",
10564=>x"002f2",
10565=>x"002f2",
10566=>x"002f2",
10567=>x"002f2",
10568=>x"002f2",
10569=>x"002f2",
10570=>x"002f3",
10571=>x"002f3",
10572=>x"002f3",
10573=>x"002f3",
10574=>x"002f3",
10575=>x"002f3",
10576=>x"002f3",
10577=>x"002f3",
10578=>x"002f3",
10579=>x"002f3",
10580=>x"002f3",
10581=>x"002f3",
10582=>x"002f3",
10583=>x"002f3",
10584=>x"002f4",
10585=>x"002f4",
10586=>x"002f4",
10587=>x"002f4",
10588=>x"002f4",
10589=>x"002f4",
10590=>x"002f4",
10591=>x"002f4",
10592=>x"002f4",
10593=>x"002f4",
10594=>x"002f4",
10595=>x"002f4",
10596=>x"002f4",
10597=>x"002f4",
10598=>x"002f5",
10599=>x"002f5",
10600=>x"002f5",
10601=>x"002f5",
10602=>x"002f5",
10603=>x"002f5",
10604=>x"002f5",
10605=>x"002f5",
10606=>x"002f5",
10607=>x"002f5",
10608=>x"002f5",
10609=>x"002f5",
10610=>x"002f5",
10611=>x"002f5",
10612=>x"002f6",
10613=>x"002f6",
10614=>x"002f6",
10615=>x"002f6",
10616=>x"002f6",
10617=>x"002f6",
10618=>x"002f6",
10619=>x"002f6",
10620=>x"002f6",
10621=>x"002f6",
10622=>x"002f6",
10623=>x"002f6",
10624=>x"002f6",
10625=>x"002f6",
10626=>x"002f7",
10627=>x"002f7",
10628=>x"002f7",
10629=>x"002f7",
10630=>x"002f7",
10631=>x"002f7",
10632=>x"002f7",
10633=>x"002f7",
10634=>x"002f7",
10635=>x"002f7",
10636=>x"002f7",
10637=>x"002f7",
10638=>x"002f7",
10639=>x"002f7",
10640=>x"002f8",
10641=>x"002f8",
10642=>x"002f8",
10643=>x"002f8",
10644=>x"002f8",
10645=>x"002f8",
10646=>x"002f8",
10647=>x"002f8",
10648=>x"002f8",
10649=>x"002f8",
10650=>x"002f8",
10651=>x"002f8",
10652=>x"002f8",
10653=>x"002f8",
10654=>x"002f9",
10655=>x"002f9",
10656=>x"002f9",
10657=>x"002f9",
10658=>x"002f9",
10659=>x"002f9",
10660=>x"002f9",
10661=>x"002f9",
10662=>x"002f9",
10663=>x"002f9",
10664=>x"002f9",
10665=>x"002f9",
10666=>x"002f9",
10667=>x"002f9",
10668=>x"002fa",
10669=>x"002fa",
10670=>x"002fa",
10671=>x"002fa",
10672=>x"002fa",
10673=>x"002fa",
10674=>x"002fa",
10675=>x"002fa",
10676=>x"002fa",
10677=>x"002fa",
10678=>x"002fa",
10679=>x"002fa",
10680=>x"002fa",
10681=>x"002fa",
10682=>x"002fb",
10683=>x"002fb",
10684=>x"002fb",
10685=>x"002fb",
10686=>x"002fb",
10687=>x"002fb",
10688=>x"002fb",
10689=>x"002fb",
10690=>x"002fb",
10691=>x"002fb",
10692=>x"002fb",
10693=>x"002fb",
10694=>x"002fb",
10695=>x"002fb",
10696=>x"002fc",
10697=>x"002fc",
10698=>x"002fc",
10699=>x"002fc",
10700=>x"002fc",
10701=>x"002fc",
10702=>x"002fc",
10703=>x"002fc",
10704=>x"002fc",
10705=>x"002fc",
10706=>x"002fc",
10707=>x"002fc",
10708=>x"002fc",
10709=>x"002fc",
10710=>x"002fd",
10711=>x"002fd",
10712=>x"002fd",
10713=>x"002fd",
10714=>x"002fd",
10715=>x"002fd",
10716=>x"002fd",
10717=>x"002fd",
10718=>x"002fd",
10719=>x"002fd",
10720=>x"002fd",
10721=>x"002fd",
10722=>x"002fd",
10723=>x"002fd",
10724=>x"002fe",
10725=>x"002fe",
10726=>x"002fe",
10727=>x"002fe",
10728=>x"002fe",
10729=>x"002fe",
10730=>x"002fe",
10731=>x"002fe",
10732=>x"002fe",
10733=>x"002fe",
10734=>x"002fe",
10735=>x"002fe",
10736=>x"002fe",
10737=>x"002fe",
10738=>x"002ff",
10739=>x"002ff",
10740=>x"002ff",
10741=>x"002ff",
10742=>x"002ff",
10743=>x"002ff",
10744=>x"002ff",
10745=>x"002ff",
10746=>x"002ff",
10747=>x"002ff",
10748=>x"002ff",
10749=>x"002ff",
10750=>x"002ff",
10751=>x"002ff",
10752=>x"00300",
10753=>x"00300",
10754=>x"00300",
10755=>x"00300",
10756=>x"00300",
10757=>x"00300",
10758=>x"00300",
10759=>x"00300",
10760=>x"00300",
10761=>x"00300",
10762=>x"00300",
10763=>x"00300",
10764=>x"00300",
10765=>x"00300",
10766=>x"00301",
10767=>x"00301",
10768=>x"00301",
10769=>x"00301",
10770=>x"00301",
10771=>x"00301",
10772=>x"00301",
10773=>x"00301",
10774=>x"00301",
10775=>x"00301",
10776=>x"00301",
10777=>x"00301",
10778=>x"00301",
10779=>x"00301",
10780=>x"00302",
10781=>x"00302",
10782=>x"00302",
10783=>x"00302",
10784=>x"00302",
10785=>x"00302",
10786=>x"00302",
10787=>x"00302",
10788=>x"00302",
10789=>x"00302",
10790=>x"00302",
10791=>x"00302",
10792=>x"00302",
10793=>x"00302",
10794=>x"00303",
10795=>x"00303",
10796=>x"00303",
10797=>x"00303",
10798=>x"00303",
10799=>x"00303",
10800=>x"00303",
10801=>x"00303",
10802=>x"00303",
10803=>x"00303",
10804=>x"00303",
10805=>x"00303",
10806=>x"00303",
10807=>x"00303",
10808=>x"00304",
10809=>x"00304",
10810=>x"00304",
10811=>x"00304",
10812=>x"00304",
10813=>x"00304",
10814=>x"00304",
10815=>x"00304",
10816=>x"00304",
10817=>x"00304",
10818=>x"00304",
10819=>x"00304",
10820=>x"00304",
10821=>x"00304",
10822=>x"00305",
10823=>x"00305",
10824=>x"00305",
10825=>x"00305",
10826=>x"00305",
10827=>x"00305",
10828=>x"00305",
10829=>x"00305",
10830=>x"00305",
10831=>x"00305",
10832=>x"00305",
10833=>x"00305",
10834=>x"00305",
10835=>x"00305",
10836=>x"00306",
10837=>x"00306",
10838=>x"00306",
10839=>x"00306",
10840=>x"00306",
10841=>x"00306",
10842=>x"00306",
10843=>x"00306",
10844=>x"00306",
10845=>x"00306",
10846=>x"00306",
10847=>x"00306",
10848=>x"00306",
10849=>x"00306",
10850=>x"00307",
10851=>x"00307",
10852=>x"00307",
10853=>x"00307",
10854=>x"00307",
10855=>x"00307",
10856=>x"00307",
10857=>x"00307",
10858=>x"00307",
10859=>x"00307",
10860=>x"00307",
10861=>x"00307",
10862=>x"00307",
10863=>x"00307",
10864=>x"00308",
10865=>x"00308",
10866=>x"00308",
10867=>x"00308",
10868=>x"00308",
10869=>x"00308",
10870=>x"00308",
10871=>x"00308",
10872=>x"00308",
10873=>x"00308",
10874=>x"00308",
10875=>x"00308",
10876=>x"00308",
10877=>x"00308",
10878=>x"00309",
10879=>x"00309",
10880=>x"00309",
10881=>x"00309",
10882=>x"00309",
10883=>x"00309",
10884=>x"00309",
10885=>x"00309",
10886=>x"00309",
10887=>x"00309",
10888=>x"00309",
10889=>x"00309",
10890=>x"00309",
10891=>x"00309",
10892=>x"0030a",
10893=>x"0030a",
10894=>x"0030a",
10895=>x"0030a",
10896=>x"0030a",
10897=>x"0030a",
10898=>x"0030a",
10899=>x"0030a",
10900=>x"0030a",
10901=>x"0030a",
10902=>x"0030a",
10903=>x"0030a",
10904=>x"0030a",
10905=>x"0030a",
10906=>x"0030b",
10907=>x"0030b",
10908=>x"0030b",
10909=>x"0030b",
10910=>x"0030b",
10911=>x"0030b",
10912=>x"0030b",
10913=>x"0030b",
10914=>x"0030b",
10915=>x"0030b",
10916=>x"0030b",
10917=>x"0030b",
10918=>x"0030b",
10919=>x"0030b",
10920=>x"0030c",
10921=>x"0030c",
10922=>x"0030c",
10923=>x"0030c",
10924=>x"0030c",
10925=>x"0030c",
10926=>x"0030c",
10927=>x"0030c",
10928=>x"0030c",
10929=>x"0030c",
10930=>x"0030c",
10931=>x"0030c",
10932=>x"0030c",
10933=>x"0030c",
10934=>x"0030d",
10935=>x"0030d",
10936=>x"0030d",
10937=>x"0030d",
10938=>x"0030d",
10939=>x"0030d",
10940=>x"0030d",
10941=>x"0030d",
10942=>x"0030d",
10943=>x"0030d",
10944=>x"0030d",
10945=>x"0030d",
10946=>x"0030d",
10947=>x"0030d",
10948=>x"0030e",
10949=>x"0030e",
10950=>x"0030e",
10951=>x"0030e",
10952=>x"0030e",
10953=>x"0030e",
10954=>x"0030e",
10955=>x"0030e",
10956=>x"0030e",
10957=>x"0030e",
10958=>x"0030e",
10959=>x"0030e",
10960=>x"0030e",
10961=>x"0030e",
10962=>x"0030f",
10963=>x"0030f",
10964=>x"0030f",
10965=>x"0030f",
10966=>x"0030f",
10967=>x"0030f",
10968=>x"0030f",
10969=>x"0030f",
10970=>x"0030f",
10971=>x"0030f",
10972=>x"0030f",
10973=>x"0030f",
10974=>x"0030f",
10975=>x"0030f",
10976=>x"00310",
10977=>x"00310",
10978=>x"00310",
10979=>x"00310",
10980=>x"00310",
10981=>x"00310",
10982=>x"00310",
10983=>x"00310",
10984=>x"00310",
10985=>x"00310",
10986=>x"00310",
10987=>x"00310",
10988=>x"00310",
10989=>x"00310",
10990=>x"00311",
10991=>x"00311",
10992=>x"00311",
10993=>x"00311",
10994=>x"00311",
10995=>x"00311",
10996=>x"00311",
10997=>x"00311",
10998=>x"00311",
10999=>x"00311",
11000=>x"00311",
11001=>x"00311",
11002=>x"00311",
11003=>x"00311",
11004=>x"00312",
11005=>x"00312",
11006=>x"00312",
11007=>x"00312",
11008=>x"00312",
11009=>x"00312",
11010=>x"00312",
11011=>x"00312",
11012=>x"00312",
11013=>x"00312",
11014=>x"00312",
11015=>x"00312",
11016=>x"00312",
11017=>x"00312",
11018=>x"00313",
11019=>x"00313",
11020=>x"00313",
11021=>x"00313",
11022=>x"00313",
11023=>x"00313",
11024=>x"00313",
11025=>x"00313",
11026=>x"00313",
11027=>x"00313",
11028=>x"00313",
11029=>x"00313",
11030=>x"00313",
11031=>x"00313",
11032=>x"00314",
11033=>x"00314",
11034=>x"00314",
11035=>x"00314",
11036=>x"00314",
11037=>x"00314",
11038=>x"00314",
11039=>x"00314",
11040=>x"00314",
11041=>x"00314",
11042=>x"00314",
11043=>x"00314",
11044=>x"00314",
11045=>x"00314",
11046=>x"00315",
11047=>x"00315",
11048=>x"00315",
11049=>x"00315",
11050=>x"00315",
11051=>x"00315",
11052=>x"00315",
11053=>x"00315",
11054=>x"00315",
11055=>x"00315",
11056=>x"00315",
11057=>x"00315",
11058=>x"00315",
11059=>x"00315",
11060=>x"00316",
11061=>x"00316",
11062=>x"00316",
11063=>x"00316",
11064=>x"00316",
11065=>x"00316",
11066=>x"00316",
11067=>x"00316",
11068=>x"00316",
11069=>x"00316",
11070=>x"00316",
11071=>x"00316",
11072=>x"00316",
11073=>x"00316",
11074=>x"00317",
11075=>x"00317",
11076=>x"00317",
11077=>x"00317",
11078=>x"00317",
11079=>x"00317",
11080=>x"00317",
11081=>x"00317",
11082=>x"00317",
11083=>x"00317",
11084=>x"00317",
11085=>x"00317",
11086=>x"00317",
11087=>x"00317",
11088=>x"00318",
11089=>x"00318",
11090=>x"00318",
11091=>x"00318",
11092=>x"00318",
11093=>x"00318",
11094=>x"00318",
11095=>x"00318",
11096=>x"00318",
11097=>x"00318",
11098=>x"00318",
11099=>x"00318",
11100=>x"00318",
11101=>x"00318",
11102=>x"00319",
11103=>x"00319",
11104=>x"00319",
11105=>x"00319",
11106=>x"00319",
11107=>x"00319",
11108=>x"00319",
11109=>x"00319",
11110=>x"00319",
11111=>x"00319",
11112=>x"00319",
11113=>x"00319",
11114=>x"00319",
11115=>x"00319",
11116=>x"0031a",
11117=>x"0031a",
11118=>x"0031a",
11119=>x"0031a",
11120=>x"0031a",
11121=>x"0031a",
11122=>x"0031a",
11123=>x"0031a",
11124=>x"0031a",
11125=>x"0031a",
11126=>x"0031a",
11127=>x"0031a",
11128=>x"0031a",
11129=>x"0031a",
11130=>x"0031b",
11131=>x"0031b",
11132=>x"0031b",
11133=>x"0031b",
11134=>x"0031b",
11135=>x"0031b",
11136=>x"0031b",
11137=>x"0031b",
11138=>x"0031b",
11139=>x"0031b",
11140=>x"0031b",
11141=>x"0031b",
11142=>x"0031b",
11143=>x"0031b",
11144=>x"0031c",
11145=>x"0031c",
11146=>x"0031c",
11147=>x"0031c",
11148=>x"0031c",
11149=>x"0031c",
11150=>x"0031c",
11151=>x"0031c",
11152=>x"0031c",
11153=>x"0031c",
11154=>x"0031c",
11155=>x"0031c",
11156=>x"0031c",
11157=>x"0031c",
11158=>x"0031d",
11159=>x"0031d",
11160=>x"0031d",
11161=>x"0031d",
11162=>x"0031d",
11163=>x"0031d",
11164=>x"0031d",
11165=>x"0031d",
11166=>x"0031d",
11167=>x"0031d",
11168=>x"0031d",
11169=>x"0031d",
11170=>x"0031d",
11171=>x"0031d",
11172=>x"0031e",
11173=>x"0031e",
11174=>x"0031e",
11175=>x"0031e",
11176=>x"0031e",
11177=>x"0031e",
11178=>x"0031e",
11179=>x"0031e",
11180=>x"0031e",
11181=>x"0031e",
11182=>x"0031e",
11183=>x"0031e",
11184=>x"0031e",
11185=>x"0031e",
11186=>x"0031f",
11187=>x"0031f",
11188=>x"0031f",
11189=>x"0031f",
11190=>x"0031f",
11191=>x"0031f",
11192=>x"0031f",
11193=>x"0031f",
11194=>x"0031f",
11195=>x"0031f",
11196=>x"0031f",
11197=>x"0031f",
11198=>x"0031f",
11199=>x"0031f",
11200=>x"00320",
11201=>x"00320",
11202=>x"00320",
11203=>x"00320",
11204=>x"00320",
11205=>x"00320",
11206=>x"00320",
11207=>x"00320",
11208=>x"00320",
11209=>x"00320",
11210=>x"00320",
11211=>x"00320",
11212=>x"00320",
11213=>x"00320",
11214=>x"00321",
11215=>x"00321",
11216=>x"00321",
11217=>x"00321",
11218=>x"00321",
11219=>x"00321",
11220=>x"00321",
11221=>x"00321",
11222=>x"00321",
11223=>x"00321",
11224=>x"00321",
11225=>x"00321",
11226=>x"00321",
11227=>x"00321",
11228=>x"00322",
11229=>x"00322",
11230=>x"00322",
11231=>x"00322",
11232=>x"00322",
11233=>x"00322",
11234=>x"00322",
11235=>x"00322",
11236=>x"00322",
11237=>x"00322",
11238=>x"00322",
11239=>x"00322",
11240=>x"00322",
11241=>x"00322",
11242=>x"00323",
11243=>x"00323",
11244=>x"00323",
11245=>x"00323",
11246=>x"00323",
11247=>x"00323",
11248=>x"00323",
11249=>x"00323",
11250=>x"00323",
11251=>x"00323",
11252=>x"00323",
11253=>x"00323",
11254=>x"00323",
11255=>x"00323",
11256=>x"00324",
11257=>x"00324",
11258=>x"00324",
11259=>x"00324",
11260=>x"00324",
11261=>x"00324",
11262=>x"00324",
11263=>x"00324",
11264=>x"00324",
11265=>x"00324",
11266=>x"00324",
11267=>x"00324",
11268=>x"00324",
11269=>x"00324",
11270=>x"00325",
11271=>x"00325",
11272=>x"00325",
11273=>x"00325",
11274=>x"00325",
11275=>x"00325",
11276=>x"00325",
11277=>x"00325",
11278=>x"00325",
11279=>x"00325",
11280=>x"00325",
11281=>x"00325",
11282=>x"00325",
11283=>x"00325",
11284=>x"00326",
11285=>x"00326",
11286=>x"00326",
11287=>x"00326",
11288=>x"00326",
11289=>x"00326",
11290=>x"00326",
11291=>x"00326",
11292=>x"00326",
11293=>x"00326",
11294=>x"00326",
11295=>x"00326",
11296=>x"00326",
11297=>x"00326",
11298=>x"00327",
11299=>x"00327",
11300=>x"00327",
11301=>x"00327",
11302=>x"00327",
11303=>x"00327",
11304=>x"00327",
11305=>x"00327",
11306=>x"00327",
11307=>x"00327",
11308=>x"00327",
11309=>x"00327",
11310=>x"00327",
11311=>x"00327",
11312=>x"00328",
11313=>x"00328",
11314=>x"00328",
11315=>x"00328",
11316=>x"00328",
11317=>x"00328",
11318=>x"00328",
11319=>x"00328",
11320=>x"00328",
11321=>x"00328",
11322=>x"00328",
11323=>x"00328",
11324=>x"00328",
11325=>x"00328",
11326=>x"00329",
11327=>x"00329",
11328=>x"00329",
11329=>x"00329",
11330=>x"00329",
11331=>x"00329",
11332=>x"00329",
11333=>x"00329",
11334=>x"00329",
11335=>x"00329",
11336=>x"00329",
11337=>x"00329",
11338=>x"00329",
11339=>x"00329",
11340=>x"0032a",
11341=>x"0032a",
11342=>x"0032a",
11343=>x"0032a",
11344=>x"0032a",
11345=>x"0032a",
11346=>x"0032a",
11347=>x"0032a",
11348=>x"0032a",
11349=>x"0032a",
11350=>x"0032a",
11351=>x"0032a",
11352=>x"0032a",
11353=>x"0032a",
11354=>x"0032b",
11355=>x"0032b",
11356=>x"0032b",
11357=>x"0032b",
11358=>x"0032b",
11359=>x"0032b",
11360=>x"0032b",
11361=>x"0032b",
11362=>x"0032b",
11363=>x"0032b",
11364=>x"0032b",
11365=>x"0032b",
11366=>x"0032b",
11367=>x"0032b",
11368=>x"0032c",
11369=>x"0032c",
11370=>x"0032c",
11371=>x"0032c",
11372=>x"0032c",
11373=>x"0032c",
11374=>x"0032c",
11375=>x"0032c",
11376=>x"0032c",
11377=>x"0032c",
11378=>x"0032c",
11379=>x"0032c",
11380=>x"0032c",
11381=>x"0032c",
11382=>x"0032d",
11383=>x"0032d",
11384=>x"0032d",
11385=>x"0032d",
11386=>x"0032d",
11387=>x"0032d",
11388=>x"0032d",
11389=>x"0032d",
11390=>x"0032d",
11391=>x"0032d",
11392=>x"0032d",
11393=>x"0032d",
11394=>x"0032d",
11395=>x"0032d",
11396=>x"0032e",
11397=>x"0032e",
11398=>x"0032e",
11399=>x"0032e",
11400=>x"0032e",
11401=>x"0032e",
11402=>x"0032e",
11403=>x"0032e",
11404=>x"0032e",
11405=>x"0032e",
11406=>x"0032e",
11407=>x"0032e",
11408=>x"0032e",
11409=>x"0032e",
11410=>x"0032f",
11411=>x"0032f",
11412=>x"0032f",
11413=>x"0032f",
11414=>x"0032f",
11415=>x"0032f",
11416=>x"0032f",
11417=>x"0032f",
11418=>x"0032f",
11419=>x"0032f",
11420=>x"0032f",
11421=>x"0032f",
11422=>x"0032f",
11423=>x"0032f",
11424=>x"00330",
11425=>x"00330",
11426=>x"00330",
11427=>x"00330",
11428=>x"00330",
11429=>x"00330",
11430=>x"00330",
11431=>x"00330",
11432=>x"00330",
11433=>x"00330",
11434=>x"00330",
11435=>x"00330",
11436=>x"00330",
11437=>x"00330",
11438=>x"00331",
11439=>x"00331",
11440=>x"00331",
11441=>x"00331",
11442=>x"00331",
11443=>x"00331",
11444=>x"00331",
11445=>x"00331",
11446=>x"00331",
11447=>x"00331",
11448=>x"00331",
11449=>x"00331",
11450=>x"00331",
11451=>x"00331",
11452=>x"00332",
11453=>x"00332",
11454=>x"00332",
11455=>x"00332",
11456=>x"00332",
11457=>x"00332",
11458=>x"00332",
11459=>x"00332",
11460=>x"00332",
11461=>x"00332",
11462=>x"00332",
11463=>x"00332",
11464=>x"00332",
11465=>x"00332",
11466=>x"00333",
11467=>x"00333",
11468=>x"00333",
11469=>x"00333",
11470=>x"00333",
11471=>x"00333",
11472=>x"00333",
11473=>x"00333",
11474=>x"00333",
11475=>x"00333",
11476=>x"00333",
11477=>x"00333",
11478=>x"00333",
11479=>x"00333",
11480=>x"00334",
11481=>x"00334",
11482=>x"00334",
11483=>x"00334",
11484=>x"00334",
11485=>x"00334",
11486=>x"00334",
11487=>x"00334",
11488=>x"00334",
11489=>x"00334",
11490=>x"00334",
11491=>x"00334",
11492=>x"00334",
11493=>x"00334",
11494=>x"00335",
11495=>x"00335",
11496=>x"00335",
11497=>x"00335",
11498=>x"00335",
11499=>x"00335",
11500=>x"00335",
11501=>x"00335",
11502=>x"00335",
11503=>x"00335",
11504=>x"00335",
11505=>x"00335",
11506=>x"00335",
11507=>x"00335",
11508=>x"00336",
11509=>x"00336",
11510=>x"00336",
11511=>x"00336",
11512=>x"00336",
11513=>x"00336",
11514=>x"00336",
11515=>x"00336",
11516=>x"00336",
11517=>x"00336",
11518=>x"00336",
11519=>x"00336",
11520=>x"00336",
11521=>x"00336",
11522=>x"00337",
11523=>x"00337",
11524=>x"00337",
11525=>x"00337",
11526=>x"00337",
11527=>x"00337",
11528=>x"00337",
11529=>x"00337",
11530=>x"00337",
11531=>x"00337",
11532=>x"00337",
11533=>x"00337",
11534=>x"00337",
11535=>x"00337",
11536=>x"00338",
11537=>x"00338",
11538=>x"00338",
11539=>x"00338",
11540=>x"00338",
11541=>x"00338",
11542=>x"00338",
11543=>x"00338",
11544=>x"00338",
11545=>x"00338",
11546=>x"00338",
11547=>x"00338",
11548=>x"00338",
11549=>x"00338",
11550=>x"00339",
11551=>x"00339",
11552=>x"00339",
11553=>x"00339",
11554=>x"00339",
11555=>x"00339",
11556=>x"00339",
11557=>x"00339",
11558=>x"00339",
11559=>x"00339",
11560=>x"00339",
11561=>x"00339",
11562=>x"00339",
11563=>x"00339",
11564=>x"0033a",
11565=>x"0033a",
11566=>x"0033a",
11567=>x"0033a",
11568=>x"0033a",
11569=>x"0033a",
11570=>x"0033a",
11571=>x"0033a",
11572=>x"0033a",
11573=>x"0033a",
11574=>x"0033a",
11575=>x"0033a",
11576=>x"0033a",
11577=>x"0033a",
11578=>x"0033b",
11579=>x"0033b",
11580=>x"0033b",
11581=>x"0033b",
11582=>x"0033b",
11583=>x"0033b",
11584=>x"0033b",
11585=>x"0033b",
11586=>x"0033b",
11587=>x"0033b",
11588=>x"0033b",
11589=>x"0033b",
11590=>x"0033b",
11591=>x"0033b",
11592=>x"0033c",
11593=>x"0033c",
11594=>x"0033c",
11595=>x"0033c",
11596=>x"0033c",
11597=>x"0033c",
11598=>x"0033c",
11599=>x"0033c",
11600=>x"0033c",
11601=>x"0033c",
11602=>x"0033c",
11603=>x"0033c",
11604=>x"0033c",
11605=>x"0033c",
11606=>x"0033d",
11607=>x"0033d",
11608=>x"0033d",
11609=>x"0033d",
11610=>x"0033d",
11611=>x"0033d",
11612=>x"0033d",
11613=>x"0033d",
11614=>x"0033d",
11615=>x"0033d",
11616=>x"0033d",
11617=>x"0033d",
11618=>x"0033d",
11619=>x"0033d",
11620=>x"0033e",
11621=>x"0033e",
11622=>x"0033e",
11623=>x"0033e",
11624=>x"0033e",
11625=>x"0033e",
11626=>x"0033e",
11627=>x"0033e",
11628=>x"0033e",
11629=>x"0033e",
11630=>x"0033e",
11631=>x"0033e",
11632=>x"0033e",
11633=>x"0033e",
11634=>x"0033f",
11635=>x"0033f",
11636=>x"0033f",
11637=>x"0033f",
11638=>x"0033f",
11639=>x"0033f",
11640=>x"0033f",
11641=>x"0033f",
11642=>x"0033f",
11643=>x"0033f",
11644=>x"0033f",
11645=>x"0033f",
11646=>x"0033f",
11647=>x"0033f",
11648=>x"00340",
11649=>x"00340",
11650=>x"00340",
11651=>x"00340",
11652=>x"00340",
11653=>x"00340",
11654=>x"00340",
11655=>x"00340",
11656=>x"00340",
11657=>x"00340",
11658=>x"00340",
11659=>x"00340",
11660=>x"00340",
11661=>x"00340",
11662=>x"00341",
11663=>x"00341",
11664=>x"00341",
11665=>x"00341",
11666=>x"00341",
11667=>x"00341",
11668=>x"00341",
11669=>x"00341",
11670=>x"00341",
11671=>x"00341",
11672=>x"00341",
11673=>x"00341",
11674=>x"00341",
11675=>x"00341",
11676=>x"00342",
11677=>x"00342",
11678=>x"00342",
11679=>x"00342",
11680=>x"00342",
11681=>x"00342",
11682=>x"00342",
11683=>x"00342",
11684=>x"00342",
11685=>x"00342",
11686=>x"00342",
11687=>x"00342",
11688=>x"00342",
11689=>x"00342",
11690=>x"00343",
11691=>x"00343",
11692=>x"00343",
11693=>x"00343",
11694=>x"00343",
11695=>x"00343",
11696=>x"00343",
11697=>x"00343",
11698=>x"00343",
11699=>x"00343",
11700=>x"00343",
11701=>x"00343",
11702=>x"00343",
11703=>x"00343",
11704=>x"00344",
11705=>x"00344",
11706=>x"00344",
11707=>x"00344",
11708=>x"00344",
11709=>x"00344",
11710=>x"00344",
11711=>x"00344",
11712=>x"00344",
11713=>x"00344",
11714=>x"00344",
11715=>x"00344",
11716=>x"00344",
11717=>x"00344",
11718=>x"00345",
11719=>x"00345",
11720=>x"00345",
11721=>x"00345",
11722=>x"00345",
11723=>x"00345",
11724=>x"00345",
11725=>x"00345",
11726=>x"00345",
11727=>x"00345",
11728=>x"00345",
11729=>x"00345",
11730=>x"00345",
11731=>x"00345",
11732=>x"00346",
11733=>x"00346",
11734=>x"00346",
11735=>x"00346",
11736=>x"00346",
11737=>x"00346",
11738=>x"00346",
11739=>x"00346",
11740=>x"00346",
11741=>x"00346",
11742=>x"00346",
11743=>x"00346",
11744=>x"00346",
11745=>x"00346",
11746=>x"00347",
11747=>x"00347",
11748=>x"00347",
11749=>x"00347",
11750=>x"00347",
11751=>x"00347",
11752=>x"00347",
11753=>x"00347",
11754=>x"00347",
11755=>x"00347",
11756=>x"00347",
11757=>x"00347",
11758=>x"00347",
11759=>x"00347",
11760=>x"00348",
11761=>x"00348",
11762=>x"00348",
11763=>x"00348",
11764=>x"00348",
11765=>x"00348",
11766=>x"00348",
11767=>x"00348",
11768=>x"00348",
11769=>x"00348",
11770=>x"00348",
11771=>x"00348",
11772=>x"00348",
11773=>x"00348",
11774=>x"00349",
11775=>x"00349",
11776=>x"00349",
11777=>x"00349",
11778=>x"00349",
11779=>x"00349",
11780=>x"00349",
11781=>x"00349",
11782=>x"00349",
11783=>x"00349",
11784=>x"00349",
11785=>x"00349",
11786=>x"00349",
11787=>x"00349",
11788=>x"0034a",
11789=>x"0034a",
11790=>x"0034a",
11791=>x"0034a",
11792=>x"0034a",
11793=>x"0034a",
11794=>x"0034a",
11795=>x"0034a",
11796=>x"0034a",
11797=>x"0034a",
11798=>x"0034a",
11799=>x"0034a",
11800=>x"0034a",
11801=>x"0034a",
11802=>x"0034b",
11803=>x"0034b",
11804=>x"0034b",
11805=>x"0034b",
11806=>x"0034b",
11807=>x"0034b",
11808=>x"0034b",
11809=>x"0034b",
11810=>x"0034b",
11811=>x"0034b",
11812=>x"0034b",
11813=>x"0034b",
11814=>x"0034b",
11815=>x"0034b",
11816=>x"0034c",
11817=>x"0034c",
11818=>x"0034c",
11819=>x"0034c",
11820=>x"0034c",
11821=>x"0034c",
11822=>x"0034c",
11823=>x"0034c",
11824=>x"0034c",
11825=>x"0034c",
11826=>x"0034c",
11827=>x"0034c",
11828=>x"0034c",
11829=>x"0034c",
11830=>x"0034d",
11831=>x"0034d",
11832=>x"0034d",
11833=>x"0034d",
11834=>x"0034d",
11835=>x"0034d",
11836=>x"0034d",
11837=>x"0034d",
11838=>x"0034d",
11839=>x"0034d",
11840=>x"0034d",
11841=>x"0034d",
11842=>x"0034d",
11843=>x"0034d",
11844=>x"0034e",
11845=>x"0034e",
11846=>x"0034e",
11847=>x"0034e",
11848=>x"0034e",
11849=>x"0034e",
11850=>x"0034e",
11851=>x"0034e",
11852=>x"0034e",
11853=>x"0034e",
11854=>x"0034e",
11855=>x"0034e",
11856=>x"0034e",
11857=>x"0034e",
11858=>x"0034f",
11859=>x"0034f",
11860=>x"0034f",
11861=>x"0034f",
11862=>x"0034f",
11863=>x"0034f",
11864=>x"0034f",
11865=>x"0034f",
11866=>x"0034f",
11867=>x"0034f",
11868=>x"0034f",
11869=>x"0034f",
11870=>x"0034f",
11871=>x"0034f",
11872=>x"00350",
11873=>x"00350",
11874=>x"00350",
11875=>x"00350",
11876=>x"00350",
11877=>x"00350",
11878=>x"00350",
11879=>x"00350",
11880=>x"00350",
11881=>x"00350",
11882=>x"00350",
11883=>x"00350",
11884=>x"00350",
11885=>x"00350",
11886=>x"00351",
11887=>x"00351",
11888=>x"00351",
11889=>x"00351",
11890=>x"00351",
11891=>x"00351",
11892=>x"00351",
11893=>x"00351",
11894=>x"00351",
11895=>x"00351",
11896=>x"00351",
11897=>x"00351",
11898=>x"00351",
11899=>x"00351",
11900=>x"00352",
11901=>x"00352",
11902=>x"00352",
11903=>x"00352",
11904=>x"00352",
11905=>x"00352",
11906=>x"00352",
11907=>x"00352",
11908=>x"00352",
11909=>x"00352",
11910=>x"00352",
11911=>x"00352",
11912=>x"00352",
11913=>x"00352",
11914=>x"00353",
11915=>x"00353",
11916=>x"00353",
11917=>x"00353",
11918=>x"00353",
11919=>x"00353",
11920=>x"00353",
11921=>x"00353",
11922=>x"00353",
11923=>x"00353",
11924=>x"00353",
11925=>x"00353",
11926=>x"00353",
11927=>x"00353",
11928=>x"00354",
11929=>x"00354",
11930=>x"00354",
11931=>x"00354",
11932=>x"00354",
11933=>x"00354",
11934=>x"00354",
11935=>x"00354",
11936=>x"00354",
11937=>x"00354",
11938=>x"00354",
11939=>x"00354",
11940=>x"00354",
11941=>x"00354",
11942=>x"00355",
11943=>x"00355",
11944=>x"00355",
11945=>x"00355",
11946=>x"00355",
11947=>x"00355",
11948=>x"00355",
11949=>x"00355",
11950=>x"00355",
11951=>x"00355",
11952=>x"00355",
11953=>x"00355",
11954=>x"00355",
11955=>x"00355",
11956=>x"00356",
11957=>x"00356",
11958=>x"00356",
11959=>x"00356",
11960=>x"00356",
11961=>x"00356",
11962=>x"00356",
11963=>x"00356",
11964=>x"00356",
11965=>x"00356",
11966=>x"00356",
11967=>x"00356",
11968=>x"00356",
11969=>x"00356",
11970=>x"00357",
11971=>x"00357",
11972=>x"00357",
11973=>x"00357",
11974=>x"00357",
11975=>x"00357",
11976=>x"00357",
11977=>x"00357",
11978=>x"00357",
11979=>x"00357",
11980=>x"00357",
11981=>x"00357",
11982=>x"00357",
11983=>x"00357",
11984=>x"00358",
11985=>x"00358",
11986=>x"00358",
11987=>x"00358",
11988=>x"00358",
11989=>x"00358",
11990=>x"00358",
11991=>x"00358",
11992=>x"00358",
11993=>x"00358",
11994=>x"00358",
11995=>x"00358",
11996=>x"00358",
11997=>x"00358",
11998=>x"00359",
11999=>x"00359",
12000=>x"00359",
12001=>x"00359",
12002=>x"00359",
12003=>x"00359",
12004=>x"00359",
12005=>x"00359",
12006=>x"00359",
12007=>x"00359",
12008=>x"00359",
12009=>x"00359",
12010=>x"00359",
12011=>x"00359",
12012=>x"0035a",
12013=>x"0035a",
12014=>x"0035a",
12015=>x"0035a",
12016=>x"0035a",
12017=>x"0035a",
12018=>x"0035a",
12019=>x"0035a",
12020=>x"0035a",
12021=>x"0035a",
12022=>x"0035a",
12023=>x"0035a",
12024=>x"0035a",
12025=>x"0035a",
12026=>x"0035b",
12027=>x"0035b",
12028=>x"0035b",
12029=>x"0035b",
12030=>x"0035b",
12031=>x"0035b",
12032=>x"0035b",
12033=>x"0035b",
12034=>x"0035b",
12035=>x"0035b",
12036=>x"0035b",
12037=>x"0035b",
12038=>x"0035b",
12039=>x"0035b",
12040=>x"0035c",
12041=>x"0035c",
12042=>x"0035c",
12043=>x"0035c",
12044=>x"0035c",
12045=>x"0035c",
12046=>x"0035c",
12047=>x"0035c",
12048=>x"0035c",
12049=>x"0035c",
12050=>x"0035c",
12051=>x"0035c",
12052=>x"0035c",
12053=>x"0035c",
12054=>x"0035d",
12055=>x"0035d",
12056=>x"0035d",
12057=>x"0035d",
12058=>x"0035d",
12059=>x"0035d",
12060=>x"0035d",
12061=>x"0035d",
12062=>x"0035d",
12063=>x"0035d",
12064=>x"0035d",
12065=>x"0035d",
12066=>x"0035d",
12067=>x"0035d",
12068=>x"0035e",
12069=>x"0035e",
12070=>x"0035e",
12071=>x"0035e",
12072=>x"0035e",
12073=>x"0035e",
12074=>x"0035e",
12075=>x"0035e",
12076=>x"0035e",
12077=>x"0035e",
12078=>x"0035e",
12079=>x"0035e",
12080=>x"0035e",
12081=>x"0035e",
12082=>x"0035f",
12083=>x"0035f",
12084=>x"0035f",
12085=>x"0035f",
12086=>x"0035f",
12087=>x"0035f",
12088=>x"0035f",
12089=>x"0035f",
12090=>x"0035f",
12091=>x"0035f",
12092=>x"0035f",
12093=>x"0035f",
12094=>x"0035f",
12095=>x"0035f",
12096=>x"00360",
12097=>x"00360",
12098=>x"00360",
12099=>x"00360",
12100=>x"00360",
12101=>x"00360",
12102=>x"00360",
12103=>x"00360",
12104=>x"00360",
12105=>x"00360",
12106=>x"00360",
12107=>x"00360",
12108=>x"00360",
12109=>x"00360",
12110=>x"00361",
12111=>x"00361",
12112=>x"00361",
12113=>x"00361",
12114=>x"00361",
12115=>x"00361",
12116=>x"00361",
12117=>x"00361",
12118=>x"00361",
12119=>x"00361",
12120=>x"00361",
12121=>x"00361",
12122=>x"00361",
12123=>x"00361",
12124=>x"00362",
12125=>x"00362",
12126=>x"00362",
12127=>x"00362",
12128=>x"00362",
12129=>x"00362",
12130=>x"00362",
12131=>x"00362",
12132=>x"00362",
12133=>x"00362",
12134=>x"00362",
12135=>x"00362",
12136=>x"00362",
12137=>x"00362",
12138=>x"00363",
12139=>x"00363",
12140=>x"00363",
12141=>x"00363",
12142=>x"00363",
12143=>x"00363",
12144=>x"00363",
12145=>x"00363",
12146=>x"00363",
12147=>x"00363",
12148=>x"00363",
12149=>x"00363",
12150=>x"00363",
12151=>x"00363",
12152=>x"00364",
12153=>x"00364",
12154=>x"00364",
12155=>x"00364",
12156=>x"00364",
12157=>x"00364",
12158=>x"00364",
12159=>x"00364",
12160=>x"00364",
12161=>x"00364",
12162=>x"00364",
12163=>x"00364",
12164=>x"00364",
12165=>x"00364",
12166=>x"00365",
12167=>x"00365",
12168=>x"00365",
12169=>x"00365",
12170=>x"00365",
12171=>x"00365",
12172=>x"00365",
12173=>x"00365",
12174=>x"00365",
12175=>x"00365",
12176=>x"00365",
12177=>x"00365",
12178=>x"00365",
12179=>x"00365",
12180=>x"00366",
12181=>x"00366",
12182=>x"00366",
12183=>x"00366",
12184=>x"00366",
12185=>x"00366",
12186=>x"00366",
12187=>x"00366",
12188=>x"00366",
12189=>x"00366",
12190=>x"00366",
12191=>x"00366",
12192=>x"00366",
12193=>x"00366",
12194=>x"00367",
12195=>x"00367",
12196=>x"00367",
12197=>x"00367",
12198=>x"00367",
12199=>x"00367",
12200=>x"00367",
12201=>x"00367",
12202=>x"00367",
12203=>x"00367",
12204=>x"00367",
12205=>x"00367",
12206=>x"00367",
12207=>x"00367",
12208=>x"00368",
12209=>x"00368",
12210=>x"00368",
12211=>x"00368",
12212=>x"00368",
12213=>x"00368",
12214=>x"00368",
12215=>x"00368",
12216=>x"00368",
12217=>x"00368",
12218=>x"00368",
12219=>x"00368",
12220=>x"00368",
12221=>x"00368",
12222=>x"00369",
12223=>x"00369",
12224=>x"00369",
12225=>x"00369",
12226=>x"00369",
12227=>x"00369",
12228=>x"00369",
12229=>x"00369",
12230=>x"00369",
12231=>x"00369",
12232=>x"00369",
12233=>x"00369",
12234=>x"00369",
12235=>x"00369",
12236=>x"0036a",
12237=>x"0036a",
12238=>x"0036a",
12239=>x"0036a",
12240=>x"0036a",
12241=>x"0036a",
12242=>x"0036a",
12243=>x"0036a",
12244=>x"0036a",
12245=>x"0036a",
12246=>x"0036a",
12247=>x"0036a",
12248=>x"0036a",
12249=>x"0036a",
12250=>x"0036b",
12251=>x"0036b",
12252=>x"0036b",
12253=>x"0036b",
12254=>x"0036b",
12255=>x"0036b",
12256=>x"0036b",
12257=>x"0036b",
12258=>x"0036b",
12259=>x"0036b",
12260=>x"0036b",
12261=>x"0036b",
12262=>x"0036b",
12263=>x"0036b",
12264=>x"0036c",
12265=>x"0036c",
12266=>x"0036c",
12267=>x"0036c",
12268=>x"0036c",
12269=>x"0036c",
12270=>x"0036c",
12271=>x"0036c",
12272=>x"0036c",
12273=>x"0036c",
12274=>x"0036c",
12275=>x"0036c",
12276=>x"0036c",
12277=>x"0036c",
12278=>x"0036d",
12279=>x"0036d",
12280=>x"0036d",
12281=>x"0036d",
12282=>x"0036d",
12283=>x"0036d",
12284=>x"0036d",
12285=>x"0036d",
12286=>x"0036d",
12287=>x"0036d",
12288=>x"0036d",
12289=>x"0036d",
12290=>x"0036d",
12291=>x"0036d",
12292=>x"0036e",
12293=>x"0036e",
12294=>x"0036e",
12295=>x"0036e",
12296=>x"0036e",
12297=>x"0036e",
12298=>x"0036e",
12299=>x"0036e",
12300=>x"0036e",
12301=>x"0036e",
12302=>x"0036e",
12303=>x"0036e",
12304=>x"0036e",
12305=>x"0036e",
12306=>x"0036f",
12307=>x"0036f",
12308=>x"0036f",
12309=>x"0036f",
12310=>x"0036f",
12311=>x"0036f",
12312=>x"0036f",
12313=>x"0036f",
12314=>x"0036f",
12315=>x"0036f",
12316=>x"0036f",
12317=>x"0036f",
12318=>x"0036f",
12319=>x"0036f",
12320=>x"00370",
12321=>x"00370",
12322=>x"00370",
12323=>x"00370",
12324=>x"00370",
12325=>x"00370",
12326=>x"00370",
12327=>x"00370",
12328=>x"00370",
12329=>x"00370",
12330=>x"00370",
12331=>x"00370",
12332=>x"00370",
12333=>x"00370",
12334=>x"00371",
12335=>x"00371",
12336=>x"00371",
12337=>x"00371",
12338=>x"00371",
12339=>x"00371",
12340=>x"00371",
12341=>x"00371",
12342=>x"00371",
12343=>x"00371",
12344=>x"00371",
12345=>x"00371",
12346=>x"00371",
12347=>x"00371",
12348=>x"00372",
12349=>x"00372",
12350=>x"00372",
12351=>x"00372",
12352=>x"00372",
12353=>x"00372",
12354=>x"00372",
12355=>x"00372",
12356=>x"00372",
12357=>x"00372",
12358=>x"00372",
12359=>x"00372",
12360=>x"00372",
12361=>x"00372",
12362=>x"00373",
12363=>x"00373",
12364=>x"00373",
12365=>x"00373",
12366=>x"00373",
12367=>x"00373",
12368=>x"00373",
12369=>x"00373",
12370=>x"00373",
12371=>x"00373",
12372=>x"00373",
12373=>x"00373",
12374=>x"00373",
12375=>x"00373",
12376=>x"00374",
12377=>x"00374",
12378=>x"00374",
12379=>x"00374",
12380=>x"00374",
12381=>x"00374",
12382=>x"00374",
12383=>x"00374",
12384=>x"00374",
12385=>x"00374",
12386=>x"00374",
12387=>x"00374",
12388=>x"00374",
12389=>x"00374",
12390=>x"00375",
12391=>x"00375",
12392=>x"00375",
12393=>x"00375",
12394=>x"00375",
12395=>x"00375",
12396=>x"00375",
12397=>x"00375",
12398=>x"00375",
12399=>x"00375",
12400=>x"00375",
12401=>x"00375",
12402=>x"00375",
12403=>x"00375",
12404=>x"00376",
12405=>x"00376",
12406=>x"00376",
12407=>x"00376",
12408=>x"00376",
12409=>x"00376",
12410=>x"00376",
12411=>x"00376",
12412=>x"00376",
12413=>x"00376",
12414=>x"00376",
12415=>x"00376",
12416=>x"00376",
12417=>x"00376",
12418=>x"00377",
12419=>x"00377",
12420=>x"00377",
12421=>x"00377",
12422=>x"00377",
12423=>x"00377",
12424=>x"00377",
12425=>x"00377",
12426=>x"00377",
12427=>x"00377",
12428=>x"00377",
12429=>x"00377",
12430=>x"00377",
12431=>x"00377",
12432=>x"00378",
12433=>x"00378",
12434=>x"00378",
12435=>x"00378",
12436=>x"00378",
12437=>x"00378",
12438=>x"00378",
12439=>x"00378",
12440=>x"00378",
12441=>x"00378",
12442=>x"00378",
12443=>x"00378",
12444=>x"00378",
12445=>x"00378",
12446=>x"00379",
12447=>x"00379",
12448=>x"00379",
12449=>x"00379",
12450=>x"00379",
12451=>x"00379",
12452=>x"00379",
12453=>x"00379",
12454=>x"00379",
12455=>x"00379",
12456=>x"00379",
12457=>x"00379",
12458=>x"00379",
12459=>x"00379",
12460=>x"0037a",
12461=>x"0037a",
12462=>x"0037a",
12463=>x"0037a",
12464=>x"0037a",
12465=>x"0037a",
12466=>x"0037a",
12467=>x"0037a",
12468=>x"0037a",
12469=>x"0037a",
12470=>x"0037a",
12471=>x"0037a",
12472=>x"0037a",
12473=>x"0037a",
12474=>x"0037b",
12475=>x"0037b",
12476=>x"0037b",
12477=>x"0037b",
12478=>x"0037b",
12479=>x"0037b",
12480=>x"0037b",
12481=>x"0037b",
12482=>x"0037b",
12483=>x"0037b",
12484=>x"0037b",
12485=>x"0037b",
12486=>x"0037b",
12487=>x"0037b",
12488=>x"0037c",
12489=>x"0037c",
12490=>x"0037c",
12491=>x"0037c",
12492=>x"0037c",
12493=>x"0037c",
12494=>x"0037c",
12495=>x"0037c",
12496=>x"0037c",
12497=>x"0037c",
12498=>x"0037c",
12499=>x"0037c",
12500=>x"0037c",
12501=>x"0037c",
12502=>x"0037d",
12503=>x"0037d",
12504=>x"0037d",
12505=>x"0037d",
12506=>x"0037d",
12507=>x"0037d",
12508=>x"0037d",
12509=>x"0037d",
12510=>x"0037d",
12511=>x"0037d",
12512=>x"0037d",
12513=>x"0037d",
12514=>x"0037d",
12515=>x"0037d",
12516=>x"0037e",
12517=>x"0037e",
12518=>x"0037e",
12519=>x"0037e",
12520=>x"0037e",
12521=>x"0037e",
12522=>x"0037e",
12523=>x"0037e",
12524=>x"0037e",
12525=>x"0037e",
12526=>x"0037e",
12527=>x"0037e",
12528=>x"0037e",
12529=>x"0037e",
12530=>x"0037f",
12531=>x"0037f",
12532=>x"0037f",
12533=>x"0037f",
12534=>x"0037f",
12535=>x"0037f",
12536=>x"0037f",
12537=>x"0037f",
12538=>x"0037f",
12539=>x"0037f",
12540=>x"0037f",
12541=>x"0037f",
12542=>x"0037f",
12543=>x"0037f",
12544=>x"00380",
12545=>x"00380",
12546=>x"00380",
12547=>x"00380",
12548=>x"00380",
12549=>x"00380",
12550=>x"00380",
12551=>x"00380",
12552=>x"00380",
12553=>x"00380",
12554=>x"00380",
12555=>x"00380",
12556=>x"00380",
12557=>x"00380",
12558=>x"00381",
12559=>x"00381",
12560=>x"00381",
12561=>x"00381",
12562=>x"00381",
12563=>x"00381",
12564=>x"00381",
12565=>x"00381",
12566=>x"00381",
12567=>x"00381",
12568=>x"00381",
12569=>x"00381",
12570=>x"00381",
12571=>x"00381",
12572=>x"00382",
12573=>x"00382",
12574=>x"00382",
12575=>x"00382",
12576=>x"00382",
12577=>x"00382",
12578=>x"00382",
12579=>x"00382",
12580=>x"00382",
12581=>x"00382",
12582=>x"00382",
12583=>x"00382",
12584=>x"00382",
12585=>x"00382",
12586=>x"00383",
12587=>x"00383",
12588=>x"00383",
12589=>x"00383",
12590=>x"00383",
12591=>x"00383",
12592=>x"00383",
12593=>x"00383",
12594=>x"00383",
12595=>x"00383",
12596=>x"00383",
12597=>x"00383",
12598=>x"00383",
12599=>x"00383",
12600=>x"00384",
12601=>x"00384",
12602=>x"00384",
12603=>x"00384",
12604=>x"00384",
12605=>x"00384",
12606=>x"00384",
12607=>x"00384",
12608=>x"00384",
12609=>x"00384",
12610=>x"00384",
12611=>x"00384",
12612=>x"00384",
12613=>x"00384",
12614=>x"00385",
12615=>x"00385",
12616=>x"00385",
12617=>x"00385",
12618=>x"00385",
12619=>x"00385",
12620=>x"00385",
12621=>x"00385",
12622=>x"00385",
12623=>x"00385",
12624=>x"00385",
12625=>x"00385",
12626=>x"00385",
12627=>x"00385",
12628=>x"00386",
12629=>x"00386",
12630=>x"00386",
12631=>x"00386",
12632=>x"00386",
12633=>x"00386",
12634=>x"00386",
12635=>x"00386",
12636=>x"00386",
12637=>x"00386",
12638=>x"00386",
12639=>x"00386",
12640=>x"00386",
12641=>x"00386",
12642=>x"00387",
12643=>x"00387",
12644=>x"00387",
12645=>x"00387",
12646=>x"00387",
12647=>x"00387",
12648=>x"00387",
12649=>x"00387",
12650=>x"00387",
12651=>x"00387",
12652=>x"00387",
12653=>x"00387",
12654=>x"00387",
12655=>x"00387",
12656=>x"00388",
12657=>x"00388",
12658=>x"00388",
12659=>x"00388",
12660=>x"00388",
12661=>x"00388",
12662=>x"00388",
12663=>x"00388",
12664=>x"00388",
12665=>x"00388",
12666=>x"00388",
12667=>x"00388",
12668=>x"00388",
12669=>x"00388",
12670=>x"00389",
12671=>x"00389",
12672=>x"00389",
12673=>x"00389",
12674=>x"00389",
12675=>x"00389",
12676=>x"00389",
12677=>x"00389",
12678=>x"00389",
12679=>x"00389",
12680=>x"00389",
12681=>x"00389",
12682=>x"00389",
12683=>x"00389",
12684=>x"0038a",
12685=>x"0038a",
12686=>x"0038a",
12687=>x"0038a",
12688=>x"0038a",
12689=>x"0038a",
12690=>x"0038a",
12691=>x"0038a",
12692=>x"0038a",
12693=>x"0038a",
12694=>x"0038a",
12695=>x"0038a",
12696=>x"0038a",
12697=>x"0038a",
12698=>x"0038b",
12699=>x"0038b",
12700=>x"0038b",
12701=>x"0038b",
12702=>x"0038b",
12703=>x"0038b",
12704=>x"0038b",
12705=>x"0038b",
12706=>x"0038b",
12707=>x"0038b",
12708=>x"0038b",
12709=>x"0038b",
12710=>x"0038b",
12711=>x"0038b",
12712=>x"0038c",
12713=>x"0038c",
12714=>x"0038c",
12715=>x"0038c",
12716=>x"0038c",
12717=>x"0038c",
12718=>x"0038c",
12719=>x"0038c",
12720=>x"0038c",
12721=>x"0038c",
12722=>x"0038c",
12723=>x"0038c",
12724=>x"0038c",
12725=>x"0038c",
12726=>x"0038d",
12727=>x"0038d",
12728=>x"0038d",
12729=>x"0038d",
12730=>x"0038d",
12731=>x"0038d",
12732=>x"0038d",
12733=>x"0038d",
12734=>x"0038d",
12735=>x"0038d",
12736=>x"0038d",
12737=>x"0038d",
12738=>x"0038d",
12739=>x"0038d",
12740=>x"0038e",
12741=>x"0038e",
12742=>x"0038e",
12743=>x"0038e",
12744=>x"0038e",
12745=>x"0038e",
12746=>x"0038e",
12747=>x"0038e",
12748=>x"0038e",
12749=>x"0038e",
12750=>x"0038e",
12751=>x"0038e",
12752=>x"0038e",
12753=>x"0038e",
12754=>x"0038f",
12755=>x"0038f",
12756=>x"0038f",
12757=>x"0038f",
12758=>x"0038f",
12759=>x"0038f",
12760=>x"0038f",
12761=>x"0038f",
12762=>x"0038f",
12763=>x"0038f",
12764=>x"0038f",
12765=>x"0038f",
12766=>x"0038f",
12767=>x"0038f",
12768=>x"00390",
12769=>x"00390",
12770=>x"00390",
12771=>x"00390",
12772=>x"00390",
12773=>x"00390",
12774=>x"00390",
12775=>x"00390",
12776=>x"00390",
12777=>x"00390",
12778=>x"00390",
12779=>x"00390",
12780=>x"00390",
12781=>x"00390",
12782=>x"00391",
12783=>x"00391",
12784=>x"00391",
12785=>x"00391",
12786=>x"00391",
12787=>x"00391",
12788=>x"00391",
12789=>x"00391",
12790=>x"00391",
12791=>x"00391",
12792=>x"00391",
12793=>x"00391",
12794=>x"00391",
12795=>x"00391",
12796=>x"00392",
12797=>x"00392",
12798=>x"00392",
12799=>x"00392",
12800=>x"00392",
12801=>x"00392",
12802=>x"00392",
12803=>x"00392",
12804=>x"00392",
12805=>x"00392",
12806=>x"00392",
12807=>x"00392",
12808=>x"00392",
12809=>x"00392",
12810=>x"00393",
12811=>x"00393",
12812=>x"00393",
12813=>x"00393",
12814=>x"00393",
12815=>x"00393",
12816=>x"00393",
12817=>x"00393",
12818=>x"00393",
12819=>x"00393",
12820=>x"00393",
12821=>x"00393",
12822=>x"00393",
12823=>x"00393",
12824=>x"00394",
12825=>x"00394",
12826=>x"00394",
12827=>x"00394",
12828=>x"00394",
12829=>x"00394",
12830=>x"00394",
12831=>x"00394",
12832=>x"00394",
12833=>x"00394",
12834=>x"00394",
12835=>x"00394",
12836=>x"00394",
12837=>x"00394",
12838=>x"00395",
12839=>x"00395",
12840=>x"00395",
12841=>x"00395",
12842=>x"00395",
12843=>x"00395",
12844=>x"00395",
12845=>x"00395",
12846=>x"00395",
12847=>x"00395",
12848=>x"00395",
12849=>x"00395",
12850=>x"00395",
12851=>x"00395",
12852=>x"00396",
12853=>x"00396",
12854=>x"00396",
12855=>x"00396",
12856=>x"00396",
12857=>x"00396",
12858=>x"00396",
12859=>x"00396",
12860=>x"00396",
12861=>x"00396",
12862=>x"00396",
12863=>x"00396",
12864=>x"00396",
12865=>x"00396",
12866=>x"00397",
12867=>x"00397",
12868=>x"00397",
12869=>x"00397",
12870=>x"00397",
12871=>x"00397",
12872=>x"00397",
12873=>x"00397",
12874=>x"00397",
12875=>x"00397",
12876=>x"00397",
12877=>x"00397",
12878=>x"00397",
12879=>x"00397",
12880=>x"00398",
12881=>x"00398",
12882=>x"00398",
12883=>x"00398",
12884=>x"00398",
12885=>x"00398",
12886=>x"00398",
12887=>x"00398",
12888=>x"00398",
12889=>x"00398",
12890=>x"00398",
12891=>x"00398",
12892=>x"00398",
12893=>x"00398",
12894=>x"00399",
12895=>x"00399",
12896=>x"00399",
12897=>x"00399",
12898=>x"00399",
12899=>x"00399",
12900=>x"00399",
12901=>x"00399",
12902=>x"00399",
12903=>x"00399",
12904=>x"00399",
12905=>x"00399",
12906=>x"00399",
12907=>x"00399",
12908=>x"0039a",
12909=>x"0039a",
12910=>x"0039a",
12911=>x"0039a",
12912=>x"0039a",
12913=>x"0039a",
12914=>x"0039a",
12915=>x"0039a",
12916=>x"0039a",
12917=>x"0039a",
12918=>x"0039a",
12919=>x"0039a",
12920=>x"0039a",
12921=>x"0039a",
12922=>x"0039b",
12923=>x"0039b",
12924=>x"0039b",
12925=>x"0039b",
12926=>x"0039b",
12927=>x"0039b",
12928=>x"0039b",
12929=>x"0039b",
12930=>x"0039b",
12931=>x"0039b",
12932=>x"0039b",
12933=>x"0039b",
12934=>x"0039b",
12935=>x"0039b",
12936=>x"0039c",
12937=>x"0039c",
12938=>x"0039c",
12939=>x"0039c",
12940=>x"0039c",
12941=>x"0039c",
12942=>x"0039c",
12943=>x"0039c",
12944=>x"0039c",
12945=>x"0039c",
12946=>x"0039c",
12947=>x"0039c",
12948=>x"0039c",
12949=>x"0039c",
12950=>x"0039d",
12951=>x"0039d",
12952=>x"0039d",
12953=>x"0039d",
12954=>x"0039d",
12955=>x"0039d",
12956=>x"0039d",
12957=>x"0039d",
12958=>x"0039d",
12959=>x"0039d",
12960=>x"0039d",
12961=>x"0039d",
12962=>x"0039d",
12963=>x"0039d",
12964=>x"0039e",
12965=>x"0039e",
12966=>x"0039e",
12967=>x"0039e",
12968=>x"0039e",
12969=>x"0039e",
12970=>x"0039e",
12971=>x"0039e",
12972=>x"0039e",
12973=>x"0039e",
12974=>x"0039e",
12975=>x"0039e",
12976=>x"0039e",
12977=>x"0039e",
12978=>x"0039f",
12979=>x"0039f",
12980=>x"0039f",
12981=>x"0039f",
12982=>x"0039f",
12983=>x"0039f",
12984=>x"0039f",
12985=>x"0039f",
12986=>x"0039f",
12987=>x"0039f",
12988=>x"0039f",
12989=>x"0039f",
12990=>x"0039f",
12991=>x"0039f",
12992=>x"003a0",
12993=>x"003a0",
12994=>x"003a0",
12995=>x"003a0",
12996=>x"003a0",
12997=>x"003a0",
12998=>x"003a0",
12999=>x"003a0",
13000=>x"003a0",
13001=>x"003a0",
13002=>x"003a0",
13003=>x"003a0",
13004=>x"003a0",
13005=>x"003a0",
13006=>x"003a1",
13007=>x"003a1",
13008=>x"003a1",
13009=>x"003a1",
13010=>x"003a1",
13011=>x"003a1",
13012=>x"003a1",
13013=>x"003a1",
13014=>x"003a1",
13015=>x"003a1",
13016=>x"003a1",
13017=>x"003a1",
13018=>x"003a1",
13019=>x"003a1",
13020=>x"003a2",
13021=>x"003a2",
13022=>x"003a2",
13023=>x"003a2",
13024=>x"003a2",
13025=>x"003a2",
13026=>x"003a2",
13027=>x"003a2",
13028=>x"003a2",
13029=>x"003a2",
13030=>x"003a2",
13031=>x"003a2",
13032=>x"003a2",
13033=>x"003a2",
13034=>x"003a3",
13035=>x"003a3",
13036=>x"003a3",
13037=>x"003a3",
13038=>x"003a3",
13039=>x"003a3",
13040=>x"003a3",
13041=>x"003a3",
13042=>x"003a3",
13043=>x"003a3",
13044=>x"003a3",
13045=>x"003a3",
13046=>x"003a3",
13047=>x"003a3",
13048=>x"003a4",
13049=>x"003a4",
13050=>x"003a4",
13051=>x"003a4",
13052=>x"003a4",
13053=>x"003a4",
13054=>x"003a4",
13055=>x"003a4",
13056=>x"003a4",
13057=>x"003a4",
13058=>x"003a4",
13059=>x"003a4",
13060=>x"003a4",
13061=>x"003a4",
13062=>x"003a5",
13063=>x"003a5",
13064=>x"003a5",
13065=>x"003a5",
13066=>x"003a5",
13067=>x"003a5",
13068=>x"003a5",
13069=>x"003a5",
13070=>x"003a5",
13071=>x"003a5",
13072=>x"003a5",
13073=>x"003a5",
13074=>x"003a5",
13075=>x"003a5",
13076=>x"003a6",
13077=>x"003a6",
13078=>x"003a6",
13079=>x"003a6",
13080=>x"003a6",
13081=>x"003a6",
13082=>x"003a6",
13083=>x"003a6",
13084=>x"003a6",
13085=>x"003a6",
13086=>x"003a6",
13087=>x"003a6",
13088=>x"003a6",
13089=>x"003a6",
13090=>x"003a7",
13091=>x"003a7",
13092=>x"003a7",
13093=>x"003a7",
13094=>x"003a7",
13095=>x"003a7",
13096=>x"003a7",
13097=>x"003a7",
13098=>x"003a7",
13099=>x"003a7",
13100=>x"003a7",
13101=>x"003a7",
13102=>x"003a7",
13103=>x"003a7",
13104=>x"003a8",
13105=>x"003a8",
13106=>x"003a8",
13107=>x"003a8",
13108=>x"003a8",
13109=>x"003a8",
13110=>x"003a8",
13111=>x"003a8",
13112=>x"003a8",
13113=>x"003a8",
13114=>x"003a8",
13115=>x"003a8",
13116=>x"003a8",
13117=>x"003a8",
13118=>x"003a9",
13119=>x"003a9",
13120=>x"003a9",
13121=>x"003a9",
13122=>x"003a9",
13123=>x"003a9",
13124=>x"003a9",
13125=>x"003a9",
13126=>x"003a9",
13127=>x"003a9",
13128=>x"003a9",
13129=>x"003a9",
13130=>x"003a9",
13131=>x"003a9",
13132=>x"003aa",
13133=>x"003aa",
13134=>x"003aa",
13135=>x"003aa",
13136=>x"003aa",
13137=>x"003aa",
13138=>x"003aa",
13139=>x"003aa",
13140=>x"003aa",
13141=>x"003aa",
13142=>x"003aa",
13143=>x"003aa",
13144=>x"003aa",
13145=>x"003aa",
13146=>x"003ab",
13147=>x"003ab",
13148=>x"003ab",
13149=>x"003ab",
13150=>x"003ab",
13151=>x"003ab",
13152=>x"003ab",
13153=>x"003ab",
13154=>x"003ab",
13155=>x"003ab",
13156=>x"003ab",
13157=>x"003ab",
13158=>x"003ab",
13159=>x"003ab",
13160=>x"003ac",
13161=>x"003ac",
13162=>x"003ac",
13163=>x"003ac",
13164=>x"003ac",
13165=>x"003ac",
13166=>x"003ac",
13167=>x"003ac",
13168=>x"003ac",
13169=>x"003ac",
13170=>x"003ac",
13171=>x"003ac",
13172=>x"003ac",
13173=>x"003ac",
13174=>x"003ad",
13175=>x"003ad",
13176=>x"003ad",
13177=>x"003ad",
13178=>x"003ad",
13179=>x"003ad",
13180=>x"003ad",
13181=>x"003ad",
13182=>x"003ad",
13183=>x"003ad",
13184=>x"003ad",
13185=>x"003ad",
13186=>x"003ad",
13187=>x"003ad",
13188=>x"003ae",
13189=>x"003ae",
13190=>x"003ae",
13191=>x"003ae",
13192=>x"003ae",
13193=>x"003ae",
13194=>x"003ae",
13195=>x"003ae",
13196=>x"003ae",
13197=>x"003ae",
13198=>x"003ae",
13199=>x"003ae",
13200=>x"003ae",
13201=>x"003ae",
13202=>x"003af",
13203=>x"003af",
13204=>x"003af",
13205=>x"003af",
13206=>x"003af",
13207=>x"003af",
13208=>x"003af",
13209=>x"003af",
13210=>x"003af",
13211=>x"003af",
13212=>x"003af",
13213=>x"003af",
13214=>x"003af",
13215=>x"003af",
13216=>x"003b0",
13217=>x"003b0",
13218=>x"003b0",
13219=>x"003b0",
13220=>x"003b0",
13221=>x"003b0",
13222=>x"003b0",
13223=>x"003b0",
13224=>x"003b0",
13225=>x"003b0",
13226=>x"003b0",
13227=>x"003b0",
13228=>x"003b0",
13229=>x"003b0",
13230=>x"003b1",
13231=>x"003b1",
13232=>x"003b1",
13233=>x"003b1",
13234=>x"003b1",
13235=>x"003b1",
13236=>x"003b1",
13237=>x"003b1",
13238=>x"003b1",
13239=>x"003b1",
13240=>x"003b1",
13241=>x"003b1",
13242=>x"003b1",
13243=>x"003b1",
13244=>x"003b2",
13245=>x"003b2",
13246=>x"003b2",
13247=>x"003b2",
13248=>x"003b2",
13249=>x"003b2",
13250=>x"003b2",
13251=>x"003b2",
13252=>x"003b2",
13253=>x"003b2",
13254=>x"003b2",
13255=>x"003b2",
13256=>x"003b2",
13257=>x"003b2",
13258=>x"003b3",
13259=>x"003b3",
13260=>x"003b3",
13261=>x"003b3",
13262=>x"003b3",
13263=>x"003b3",
13264=>x"003b3",
13265=>x"003b3",
13266=>x"003b3",
13267=>x"003b3",
13268=>x"003b3",
13269=>x"003b3",
13270=>x"003b3",
13271=>x"003b3",
13272=>x"003b4",
13273=>x"003b4",
13274=>x"003b4",
13275=>x"003b4",
13276=>x"003b4",
13277=>x"003b4",
13278=>x"003b4",
13279=>x"003b4",
13280=>x"003b4",
13281=>x"003b4",
13282=>x"003b4",
13283=>x"003b4",
13284=>x"003b4",
13285=>x"003b4",
13286=>x"003b5",
13287=>x"003b5",
13288=>x"003b5",
13289=>x"003b5",
13290=>x"003b5",
13291=>x"003b5",
13292=>x"003b5",
13293=>x"003b5",
13294=>x"003b5",
13295=>x"003b5",
13296=>x"003b5",
13297=>x"003b5",
13298=>x"003b5",
13299=>x"003b5",
13300=>x"003b6",
13301=>x"003b6",
13302=>x"003b6",
13303=>x"003b6",
13304=>x"003b6",
13305=>x"003b6",
13306=>x"003b6",
13307=>x"003b6",
13308=>x"003b6",
13309=>x"003b6",
13310=>x"003b6",
13311=>x"003b6",
13312=>x"003b6",
13313=>x"003b6",
13314=>x"003b7",
13315=>x"003b7",
13316=>x"003b7",
13317=>x"003b7",
13318=>x"003b7",
13319=>x"003b7",
13320=>x"003b7",
13321=>x"003b7",
13322=>x"003b7",
13323=>x"003b7",
13324=>x"003b7",
13325=>x"003b7",
13326=>x"003b7",
13327=>x"003b7",
13328=>x"003b8",
13329=>x"003b8",
13330=>x"003b8",
13331=>x"003b8",
13332=>x"003b8",
13333=>x"003b8",
13334=>x"003b8",
13335=>x"003b8",
13336=>x"003b8",
13337=>x"003b8",
13338=>x"003b8",
13339=>x"003b8",
13340=>x"003b8",
13341=>x"003b8",
13342=>x"003b9",
13343=>x"003b9",
13344=>x"003b9",
13345=>x"003b9",
13346=>x"003b9",
13347=>x"003b9",
13348=>x"003b9",
13349=>x"003b9",
13350=>x"003b9",
13351=>x"003b9",
13352=>x"003b9",
13353=>x"003b9",
13354=>x"003b9",
13355=>x"003b9",
13356=>x"003ba",
13357=>x"003ba",
13358=>x"003ba",
13359=>x"003ba",
13360=>x"003ba",
13361=>x"003ba",
13362=>x"003ba",
13363=>x"003ba",
13364=>x"003ba",
13365=>x"003ba",
13366=>x"003ba",
13367=>x"003ba",
13368=>x"003ba",
13369=>x"003ba",
13370=>x"003bb",
13371=>x"003bb",
13372=>x"003bb",
13373=>x"003bb",
13374=>x"003bb",
13375=>x"003bb",
13376=>x"003bb",
13377=>x"003bb",
13378=>x"003bb",
13379=>x"003bb",
13380=>x"003bb",
13381=>x"003bb",
13382=>x"003bb",
13383=>x"003bb",
13384=>x"003bc",
13385=>x"003bc",
13386=>x"003bc",
13387=>x"003bc",
13388=>x"003bc",
13389=>x"003bc",
13390=>x"003bc",
13391=>x"003bc",
13392=>x"003bc",
13393=>x"003bc",
13394=>x"003bc",
13395=>x"003bc",
13396=>x"003bc",
13397=>x"003bc",
13398=>x"003bd",
13399=>x"003bd",
13400=>x"003bd",
13401=>x"003bd",
13402=>x"003bd",
13403=>x"003bd",
13404=>x"003bd",
13405=>x"003bd",
13406=>x"003bd",
13407=>x"003bd",
13408=>x"003bd",
13409=>x"003bd",
13410=>x"003bd",
13411=>x"003bd",
13412=>x"003be",
13413=>x"003be",
13414=>x"003be",
13415=>x"003be",
13416=>x"003be",
13417=>x"003be",
13418=>x"003be",
13419=>x"003be",
13420=>x"003be",
13421=>x"003be",
13422=>x"003be",
13423=>x"003be",
13424=>x"003be",
13425=>x"003be",
13426=>x"003bf",
13427=>x"003bf",
13428=>x"003bf",
13429=>x"003bf",
13430=>x"003bf",
13431=>x"003bf",
13432=>x"003bf",
13433=>x"003bf",
13434=>x"003bf",
13435=>x"003bf",
13436=>x"003bf",
13437=>x"003bf",
13438=>x"003bf",
13439=>x"003bf",
13440=>x"003c0",
13441=>x"003c0",
13442=>x"003c0",
13443=>x"003c0",
13444=>x"003c0",
13445=>x"003c0",
13446=>x"003c0",
13447=>x"003c0",
13448=>x"003c0",
13449=>x"003c0",
13450=>x"003c0",
13451=>x"003c0",
13452=>x"003c0",
13453=>x"003c0",
13454=>x"003c1",
13455=>x"003c1",
13456=>x"003c1",
13457=>x"003c1",
13458=>x"003c1",
13459=>x"003c1",
13460=>x"003c1",
13461=>x"003c1",
13462=>x"003c1",
13463=>x"003c1",
13464=>x"003c1",
13465=>x"003c1",
13466=>x"003c1",
13467=>x"003c1",
13468=>x"003c2",
13469=>x"003c2",
13470=>x"003c2",
13471=>x"003c2",
13472=>x"003c2",
13473=>x"003c2",
13474=>x"003c2",
13475=>x"003c2",
13476=>x"003c2",
13477=>x"003c2",
13478=>x"003c2",
13479=>x"003c2",
13480=>x"003c2",
13481=>x"003c2",
13482=>x"003c3",
13483=>x"003c3",
13484=>x"003c3",
13485=>x"003c3",
13486=>x"003c3",
13487=>x"003c3",
13488=>x"003c3",
13489=>x"003c3",
13490=>x"003c3",
13491=>x"003c3",
13492=>x"003c3",
13493=>x"003c3",
13494=>x"003c3",
13495=>x"003c3",
13496=>x"003c4",
13497=>x"003c4",
13498=>x"003c4",
13499=>x"003c4",
13500=>x"003c4",
13501=>x"003c4",
13502=>x"003c4",
13503=>x"003c4",
13504=>x"003c4",
13505=>x"003c4",
13506=>x"003c4",
13507=>x"003c4",
13508=>x"003c4",
13509=>x"003c4",
13510=>x"003c5",
13511=>x"003c5",
13512=>x"003c5",
13513=>x"003c5",
13514=>x"003c5",
13515=>x"003c5",
13516=>x"003c5",
13517=>x"003c5",
13518=>x"003c5",
13519=>x"003c5",
13520=>x"003c5",
13521=>x"003c5",
13522=>x"003c5",
13523=>x"003c5",
13524=>x"003c6",
13525=>x"003c6",
13526=>x"003c6",
13527=>x"003c6",
13528=>x"003c6",
13529=>x"003c6",
13530=>x"003c6",
13531=>x"003c6",
13532=>x"003c6",
13533=>x"003c6",
13534=>x"003c6",
13535=>x"003c6",
13536=>x"003c6",
13537=>x"003c6",
13538=>x"003c7",
13539=>x"003c7",
13540=>x"003c7",
13541=>x"003c7",
13542=>x"003c7",
13543=>x"003c7",
13544=>x"003c7",
13545=>x"003c7",
13546=>x"003c7",
13547=>x"003c7",
13548=>x"003c7",
13549=>x"003c7",
13550=>x"003c7",
13551=>x"003c7",
13552=>x"003c8",
13553=>x"003c8",
13554=>x"003c8",
13555=>x"003c8",
13556=>x"003c8",
13557=>x"003c8",
13558=>x"003c8",
13559=>x"003c8",
13560=>x"003c8",
13561=>x"003c8",
13562=>x"003c8",
13563=>x"003c8",
13564=>x"003c8",
13565=>x"003c8",
13566=>x"003c9",
13567=>x"003c9",
13568=>x"003c9",
13569=>x"003c9",
13570=>x"003c9",
13571=>x"003c9",
13572=>x"003c9",
13573=>x"003c9",
13574=>x"003c9",
13575=>x"003c9",
13576=>x"003c9",
13577=>x"003c9",
13578=>x"003c9",
13579=>x"003c9",
13580=>x"003ca",
13581=>x"003ca",
13582=>x"003ca",
13583=>x"003ca",
13584=>x"003ca",
13585=>x"003ca",
13586=>x"003ca",
13587=>x"003ca",
13588=>x"003ca",
13589=>x"003ca",
13590=>x"003ca",
13591=>x"003ca",
13592=>x"003ca",
13593=>x"003ca",
13594=>x"003cb",
13595=>x"003cb",
13596=>x"003cb",
13597=>x"003cb",
13598=>x"003cb",
13599=>x"003cb",
13600=>x"003cb",
13601=>x"003cb",
13602=>x"003cb",
13603=>x"003cb",
13604=>x"003cb",
13605=>x"003cb",
13606=>x"003cb",
13607=>x"003cb",
13608=>x"003cc",
13609=>x"003cc",
13610=>x"003cc",
13611=>x"003cc",
13612=>x"003cc",
13613=>x"003cc",
13614=>x"003cc",
13615=>x"003cc",
13616=>x"003cc",
13617=>x"003cc",
13618=>x"003cc",
13619=>x"003cc",
13620=>x"003cc",
13621=>x"003cc",
13622=>x"003cd",
13623=>x"003cd",
13624=>x"003cd",
13625=>x"003cd",
13626=>x"003cd",
13627=>x"003cd",
13628=>x"003cd",
13629=>x"003cd",
13630=>x"003cd",
13631=>x"003cd",
13632=>x"003cd",
13633=>x"003cd",
13634=>x"003cd",
13635=>x"003cd",
13636=>x"003ce",
13637=>x"003ce",
13638=>x"003ce",
13639=>x"003ce",
13640=>x"003ce",
13641=>x"003ce",
13642=>x"003ce",
13643=>x"003ce",
13644=>x"003ce",
13645=>x"003ce",
13646=>x"003ce",
13647=>x"003ce",
13648=>x"003ce",
13649=>x"003ce",
13650=>x"003cf",
13651=>x"003cf",
13652=>x"003cf",
13653=>x"003cf",
13654=>x"003cf",
13655=>x"003cf",
13656=>x"003cf",
13657=>x"003cf",
13658=>x"003cf",
13659=>x"003cf",
13660=>x"003cf",
13661=>x"003cf",
13662=>x"003cf",
13663=>x"003cf",
13664=>x"003d0",
13665=>x"003d0",
13666=>x"003d0",
13667=>x"003d0",
13668=>x"003d0",
13669=>x"003d0",
13670=>x"003d0",
13671=>x"003d0",
13672=>x"003d0",
13673=>x"003d0",
13674=>x"003d0",
13675=>x"003d0",
13676=>x"003d0",
13677=>x"003d0",
13678=>x"003d1",
13679=>x"003d1",
13680=>x"003d1",
13681=>x"003d1",
13682=>x"003d1",
13683=>x"003d1",
13684=>x"003d1",
13685=>x"003d1",
13686=>x"003d1",
13687=>x"003d1",
13688=>x"003d1",
13689=>x"003d1",
13690=>x"003d1",
13691=>x"003d1",
13692=>x"003d2",
13693=>x"003d2",
13694=>x"003d2",
13695=>x"003d2",
13696=>x"003d2",
13697=>x"003d2",
13698=>x"003d2",
13699=>x"003d2",
13700=>x"003d2",
13701=>x"003d2",
13702=>x"003d2",
13703=>x"003d2",
13704=>x"003d2",
13705=>x"003d2",
13706=>x"003d3",
13707=>x"003d3",
13708=>x"003d3",
13709=>x"003d3",
13710=>x"003d3",
13711=>x"003d3",
13712=>x"003d3",
13713=>x"003d3",
13714=>x"003d3",
13715=>x"003d3",
13716=>x"003d3",
13717=>x"003d3",
13718=>x"003d3",
13719=>x"003d3",
13720=>x"003d4",
13721=>x"003d4",
13722=>x"003d4",
13723=>x"003d4",
13724=>x"003d4",
13725=>x"003d4",
13726=>x"003d4",
13727=>x"003d4",
13728=>x"003d4",
13729=>x"003d4",
13730=>x"003d4",
13731=>x"003d4",
13732=>x"003d4",
13733=>x"003d4",
13734=>x"003d5",
13735=>x"003d5",
13736=>x"003d5",
13737=>x"003d5",
13738=>x"003d5",
13739=>x"003d5",
13740=>x"003d5",
13741=>x"003d5",
13742=>x"003d5",
13743=>x"003d5",
13744=>x"003d5",
13745=>x"003d5",
13746=>x"003d5",
13747=>x"003d5",
13748=>x"003d6",
13749=>x"003d6",
13750=>x"003d6",
13751=>x"003d6",
13752=>x"003d6",
13753=>x"003d6",
13754=>x"003d6",
13755=>x"003d6",
13756=>x"003d6",
13757=>x"003d6",
13758=>x"003d6",
13759=>x"003d6",
13760=>x"003d6",
13761=>x"003d6",
13762=>x"003d7",
13763=>x"003d7",
13764=>x"003d7",
13765=>x"003d7",
13766=>x"003d7",
13767=>x"003d7",
13768=>x"003d7",
13769=>x"003d7",
13770=>x"003d7",
13771=>x"003d7",
13772=>x"003d7",
13773=>x"003d7",
13774=>x"003d7",
13775=>x"003d7",
13776=>x"003d8",
13777=>x"003d8",
13778=>x"003d8",
13779=>x"003d8",
13780=>x"003d8",
13781=>x"003d8",
13782=>x"003d8",
13783=>x"003d8",
13784=>x"003d8",
13785=>x"003d8",
13786=>x"003d8",
13787=>x"003d8",
13788=>x"003d8",
13789=>x"003d8",
13790=>x"003d9",
13791=>x"003d9",
13792=>x"003d9",
13793=>x"003d9",
13794=>x"003d9",
13795=>x"003d9",
13796=>x"003d9",
13797=>x"003d9",
13798=>x"003d9",
13799=>x"003d9",
13800=>x"003d9",
13801=>x"003d9",
13802=>x"003d9",
13803=>x"003d9",
13804=>x"003da",
13805=>x"003da",
13806=>x"003da",
13807=>x"003da",
13808=>x"003da",
13809=>x"003da",
13810=>x"003da",
13811=>x"003da",
13812=>x"003da",
13813=>x"003da",
13814=>x"003da",
13815=>x"003da",
13816=>x"003da",
13817=>x"003da",
13818=>x"003db",
13819=>x"003db",
13820=>x"003db",
13821=>x"003db",
13822=>x"003db",
13823=>x"003db",
13824=>x"003db",
13825=>x"003db",
13826=>x"003db",
13827=>x"003db",
13828=>x"003db",
13829=>x"003db",
13830=>x"003db",
13831=>x"003db",
13832=>x"003dc",
13833=>x"003dc",
13834=>x"003dc",
13835=>x"003dc",
13836=>x"003dc",
13837=>x"003dc",
13838=>x"003dc",
13839=>x"003dc",
13840=>x"003dc",
13841=>x"003dc",
13842=>x"003dc",
13843=>x"003dc",
13844=>x"003dc",
13845=>x"003dc",
13846=>x"003dd",
13847=>x"003dd",
13848=>x"003dd",
13849=>x"003dd",
13850=>x"003dd",
13851=>x"003dd",
13852=>x"003dd",
13853=>x"003dd",
13854=>x"003dd",
13855=>x"003dd",
13856=>x"003dd",
13857=>x"003dd",
13858=>x"003dd",
13859=>x"003dd",
13860=>x"003de",
13861=>x"003de",
13862=>x"003de",
13863=>x"003de",
13864=>x"003de",
13865=>x"003de",
13866=>x"003de",
13867=>x"003de",
13868=>x"003de",
13869=>x"003de",
13870=>x"003de",
13871=>x"003de",
13872=>x"003de",
13873=>x"003de",
13874=>x"003df",
13875=>x"003df",
13876=>x"003df",
13877=>x"003df",
13878=>x"003df",
13879=>x"003df",
13880=>x"003df",
13881=>x"003df",
13882=>x"003df",
13883=>x"003df",
13884=>x"003df",
13885=>x"003df",
13886=>x"003df",
13887=>x"003df",
13888=>x"003e0",
13889=>x"003e0",
13890=>x"003e0",
13891=>x"003e0",
13892=>x"003e0",
13893=>x"003e0",
13894=>x"003e0",
13895=>x"003e0",
13896=>x"003e0",
13897=>x"003e0",
13898=>x"003e0",
13899=>x"003e0",
13900=>x"003e0",
13901=>x"003e0",
13902=>x"003e1",
13903=>x"003e1",
13904=>x"003e1",
13905=>x"003e1",
13906=>x"003e1",
13907=>x"003e1",
13908=>x"003e1",
13909=>x"003e1",
13910=>x"003e1",
13911=>x"003e1",
13912=>x"003e1",
13913=>x"003e1",
13914=>x"003e1",
13915=>x"003e1",
13916=>x"003e2",
13917=>x"003e2",
13918=>x"003e2",
13919=>x"003e2",
13920=>x"003e2",
13921=>x"003e2",
13922=>x"003e2",
13923=>x"003e2",
13924=>x"003e2",
13925=>x"003e2",
13926=>x"003e2",
13927=>x"003e2",
13928=>x"003e2",
13929=>x"003e2",
13930=>x"003e3",
13931=>x"003e3",
13932=>x"003e3",
13933=>x"003e3",
13934=>x"003e3",
13935=>x"003e3",
13936=>x"003e3",
13937=>x"003e3",
13938=>x"003e3",
13939=>x"003e3",
13940=>x"003e3",
13941=>x"003e3",
13942=>x"003e3",
13943=>x"003e3",
13944=>x"003e4",
13945=>x"003e4",
13946=>x"003e4",
13947=>x"003e4",
13948=>x"003e4",
13949=>x"003e4",
13950=>x"003e4",
13951=>x"003e4",
13952=>x"003e4",
13953=>x"003e4",
13954=>x"003e4",
13955=>x"003e4",
13956=>x"003e4",
13957=>x"003e4",
13958=>x"003e5",
13959=>x"003e5",
13960=>x"003e5",
13961=>x"003e5",
13962=>x"003e5",
13963=>x"003e5",
13964=>x"003e5",
13965=>x"003e5",
13966=>x"003e5",
13967=>x"003e5",
13968=>x"003e5",
13969=>x"003e5",
13970=>x"003e5",
13971=>x"003e5",
13972=>x"003e6",
13973=>x"003e6",
13974=>x"003e6",
13975=>x"003e6",
13976=>x"003e6",
13977=>x"003e6",
13978=>x"003e6",
13979=>x"003e6",
13980=>x"003e6",
13981=>x"003e6",
13982=>x"003e6",
13983=>x"003e6",
13984=>x"003e6",
13985=>x"003e6",
13986=>x"003e7",
13987=>x"003e7",
13988=>x"003e7",
13989=>x"003e7",
13990=>x"003e7",
13991=>x"003e7",
13992=>x"003e7",
13993=>x"003e7",
13994=>x"003e7",
13995=>x"003e7",
13996=>x"003e7",
13997=>x"003e7",
13998=>x"003e7",
13999=>x"003e7",
14000=>x"003e8",
14001=>x"003e8",
14002=>x"003e8",
14003=>x"003e8",
14004=>x"003e8",
14005=>x"003e8",
14006=>x"003e8",
14007=>x"003e8",
14008=>x"003e8",
14009=>x"003e8",
14010=>x"003e8",
14011=>x"003e8",
14012=>x"003e8",
14013=>x"003e8",
14014=>x"003e9",
14015=>x"003e9",
14016=>x"003e9",
14017=>x"003e9",
14018=>x"003e9",
14019=>x"003e9",
14020=>x"003e9",
14021=>x"003e9",
14022=>x"003e9",
14023=>x"003e9",
14024=>x"003e9",
14025=>x"003e9",
14026=>x"003e9",
14027=>x"003e9",
14028=>x"003ea",
14029=>x"003ea",
14030=>x"003ea",
14031=>x"003ea",
14032=>x"003ea",
14033=>x"003ea",
14034=>x"003ea",
14035=>x"003ea",
14036=>x"003ea",
14037=>x"003ea",
14038=>x"003ea",
14039=>x"003ea",
14040=>x"003ea",
14041=>x"003ea",
14042=>x"003eb",
14043=>x"003eb",
14044=>x"003eb",
14045=>x"003eb",
14046=>x"003eb",
14047=>x"003eb",
14048=>x"003eb",
14049=>x"003eb",
14050=>x"003eb",
14051=>x"003eb",
14052=>x"003eb",
14053=>x"003eb",
14054=>x"003eb",
14055=>x"003eb",
14056=>x"003ec",
14057=>x"003ec",
14058=>x"003ec",
14059=>x"003ec",
14060=>x"003ec",
14061=>x"003ec",
14062=>x"003ec",
14063=>x"003ec",
14064=>x"003ec",
14065=>x"003ec",
14066=>x"003ec",
14067=>x"003ec",
14068=>x"003ec",
14069=>x"003ec",
14070=>x"003ed",
14071=>x"003ed",
14072=>x"003ed",
14073=>x"003ed",
14074=>x"003ed",
14075=>x"003ed",
14076=>x"003ed",
14077=>x"003ed",
14078=>x"003ed",
14079=>x"003ed",
14080=>x"003ed",
14081=>x"003ed",
14082=>x"003ed",
14083=>x"003ed",
14084=>x"003ee",
14085=>x"003ee",
14086=>x"003ee",
14087=>x"003ee",
14088=>x"003ee",
14089=>x"003ee",
14090=>x"003ee",
14091=>x"003ee",
14092=>x"003ee",
14093=>x"003ee",
14094=>x"003ee",
14095=>x"003ee",
14096=>x"003ee",
14097=>x"003ee",
14098=>x"003ef",
14099=>x"003ef",
14100=>x"003ef",
14101=>x"003ef",
14102=>x"003ef",
14103=>x"003ef",
14104=>x"003ef",
14105=>x"003ef",
14106=>x"003ef",
14107=>x"003ef",
14108=>x"003ef",
14109=>x"003ef",
14110=>x"003ef",
14111=>x"003ef",
14112=>x"003f0",
14113=>x"003f0",
14114=>x"003f0",
14115=>x"003f0",
14116=>x"003f0",
14117=>x"003f0",
14118=>x"003f0",
14119=>x"003f0",
14120=>x"003f0",
14121=>x"003f0",
14122=>x"003f0",
14123=>x"003f0",
14124=>x"003f0",
14125=>x"003f0",
14126=>x"003f1",
14127=>x"003f1",
14128=>x"003f1",
14129=>x"003f1",
14130=>x"003f1",
14131=>x"003f1",
14132=>x"003f1",
14133=>x"003f1",
14134=>x"003f1",
14135=>x"003f1",
14136=>x"003f1",
14137=>x"003f1",
14138=>x"003f1",
14139=>x"003f1",
14140=>x"003f2",
14141=>x"003f2",
14142=>x"003f2",
14143=>x"003f2",
14144=>x"003f2",
14145=>x"003f2",
14146=>x"003f2",
14147=>x"003f2",
14148=>x"003f2",
14149=>x"003f2",
14150=>x"003f2",
14151=>x"003f2",
14152=>x"003f2",
14153=>x"003f2",
14154=>x"003f3",
14155=>x"003f3",
14156=>x"003f3",
14157=>x"003f3",
14158=>x"003f3",
14159=>x"003f3",
14160=>x"003f3",
14161=>x"003f3",
14162=>x"003f3",
14163=>x"003f3",
14164=>x"003f3",
14165=>x"003f3",
14166=>x"003f3",
14167=>x"003f3",
14168=>x"003f4",
14169=>x"003f4",
14170=>x"003f4",
14171=>x"003f4",
14172=>x"003f4",
14173=>x"003f4",
14174=>x"003f4",
14175=>x"003f4",
14176=>x"003f4",
14177=>x"003f4",
14178=>x"003f4",
14179=>x"003f4",
14180=>x"003f4",
14181=>x"003f4",
14182=>x"003f5",
14183=>x"003f5",
14184=>x"003f5",
14185=>x"003f5",
14186=>x"003f5",
14187=>x"003f5",
14188=>x"003f5",
14189=>x"003f5",
14190=>x"003f5",
14191=>x"003f5",
14192=>x"003f5",
14193=>x"003f5",
14194=>x"003f5",
14195=>x"003f5",
14196=>x"003f6",
14197=>x"003f6",
14198=>x"003f6",
14199=>x"003f6",
14200=>x"003f6",
14201=>x"003f6",
14202=>x"003f6",
14203=>x"003f6",
14204=>x"003f6",
14205=>x"003f6",
14206=>x"003f6",
14207=>x"003f6",
14208=>x"003f6",
14209=>x"003f6",
14210=>x"003f7",
14211=>x"003f7",
14212=>x"003f7",
14213=>x"003f7",
14214=>x"003f7",
14215=>x"003f7",
14216=>x"003f7",
14217=>x"003f7",
14218=>x"003f7",
14219=>x"003f7",
14220=>x"003f7",
14221=>x"003f7",
14222=>x"003f7",
14223=>x"003f7",
14224=>x"003f8",
14225=>x"003f8",
14226=>x"003f8",
14227=>x"003f8",
14228=>x"003f8",
14229=>x"003f8",
14230=>x"003f8",
14231=>x"003f8",
14232=>x"003f8",
14233=>x"003f8",
14234=>x"003f8",
14235=>x"003f8",
14236=>x"003f8",
14237=>x"003f8",
14238=>x"003f9",
14239=>x"003f9",
14240=>x"003f9",
14241=>x"003f9",
14242=>x"003f9",
14243=>x"003f9",
14244=>x"003f9",
14245=>x"003f9",
14246=>x"003f9",
14247=>x"003f9",
14248=>x"003f9",
14249=>x"003f9",
14250=>x"003f9",
14251=>x"003f9",
14252=>x"003fa",
14253=>x"003fa",
14254=>x"003fa",
14255=>x"003fa",
14256=>x"003fa",
14257=>x"003fa",
14258=>x"003fa",
14259=>x"003fa",
14260=>x"003fa",
14261=>x"003fa",
14262=>x"003fa",
14263=>x"003fa",
14264=>x"003fa",
14265=>x"003fa",
14266=>x"003fb",
14267=>x"003fb",
14268=>x"003fb",
14269=>x"003fb",
14270=>x"003fb",
14271=>x"003fb",
14272=>x"003fb",
14273=>x"003fb",
14274=>x"003fb",
14275=>x"003fb",
14276=>x"003fb",
14277=>x"003fb",
14278=>x"003fb",
14279=>x"003fb",
14280=>x"003fc",
14281=>x"003fc",
14282=>x"003fc",
14283=>x"003fc",
14284=>x"003fc",
14285=>x"003fc",
14286=>x"003fc",
14287=>x"003fc",
14288=>x"003fc",
14289=>x"003fc",
14290=>x"003fc",
14291=>x"003fc",
14292=>x"003fc",
14293=>x"003fc",
14294=>x"003fd",
14295=>x"003fd",
14296=>x"003fd",
14297=>x"003fd",
14298=>x"003fd",
14299=>x"003fd",
14300=>x"003fd",
14301=>x"003fd",
14302=>x"003fd",
14303=>x"003fd",
14304=>x"003fd",
14305=>x"003fd",
14306=>x"003fd",
14307=>x"003fd",
14308=>x"003fe",
14309=>x"003fe",
14310=>x"003fe",
14311=>x"003fe",
14312=>x"003fe",
14313=>x"003fe",
14314=>x"003fe",
14315=>x"003fe",
14316=>x"003fe",
14317=>x"003fe",
14318=>x"003fe",
14319=>x"003fe",
14320=>x"003fe",
14321=>x"003fe",
14322=>x"003ff",
14323=>x"003ff",
14324=>x"003ff",
14325=>x"003ff",
14326=>x"003ff",
14327=>x"003ff",
14328=>x"003ff",
14329=>x"003ff",
14330=>x"003ff",
14331=>x"003ff",
14332=>x"003ff",
14333=>x"003ff",
14334=>x"003ff",
14335=>x"003ff",
14336=>x"00400",
14337=>x"00400",
14338=>x"00400",
14339=>x"00400",
14340=>x"00400",
14341=>x"00400",
14342=>x"00400",
14343=>x"00400",
14344=>x"00400",
14345=>x"00400",
14346=>x"00400",
14347=>x"00400",
14348=>x"00400",
14349=>x"00400",
14350=>x"00401",
14351=>x"00401",
14352=>x"00401",
14353=>x"00401",
14354=>x"00401",
14355=>x"00401",
14356=>x"00401",
14357=>x"00401",
14358=>x"00401",
14359=>x"00401",
14360=>x"00401",
14361=>x"00401",
14362=>x"00401",
14363=>x"00401",
14364=>x"00402",
14365=>x"00402",
14366=>x"00402",
14367=>x"00402",
14368=>x"00402",
14369=>x"00402",
14370=>x"00402",
14371=>x"00402",
14372=>x"00402",
14373=>x"00402",
14374=>x"00402",
14375=>x"00402",
14376=>x"00402",
14377=>x"00402",
14378=>x"00403",
14379=>x"00403",
14380=>x"00403",
14381=>x"00403",
14382=>x"00403",
14383=>x"00403",
14384=>x"00403",
14385=>x"00403",
14386=>x"00403",
14387=>x"00403",
14388=>x"00403",
14389=>x"00403",
14390=>x"00403",
14391=>x"00403",
14392=>x"00404",
14393=>x"00404",
14394=>x"00404",
14395=>x"00404",
14396=>x"00404",
14397=>x"00404",
14398=>x"00404",
14399=>x"00404",
14400=>x"00404",
14401=>x"00404",
14402=>x"00404",
14403=>x"00404",
14404=>x"00404",
14405=>x"00404",
14406=>x"00405",
14407=>x"00405",
14408=>x"00405",
14409=>x"00405",
14410=>x"00405",
14411=>x"00405",
14412=>x"00405",
14413=>x"00405",
14414=>x"00405",
14415=>x"00405",
14416=>x"00405",
14417=>x"00405",
14418=>x"00405",
14419=>x"00405",
14420=>x"00406",
14421=>x"00406",
14422=>x"00406",
14423=>x"00406",
14424=>x"00406",
14425=>x"00406",
14426=>x"00406",
14427=>x"00406",
14428=>x"00406",
14429=>x"00406",
14430=>x"00406",
14431=>x"00406",
14432=>x"00406",
14433=>x"00406",
14434=>x"00407",
14435=>x"00407",
14436=>x"00407",
14437=>x"00407",
14438=>x"00407",
14439=>x"00407",
14440=>x"00407",
14441=>x"00407",
14442=>x"00407",
14443=>x"00407",
14444=>x"00407",
14445=>x"00407",
14446=>x"00407",
14447=>x"00407",
14448=>x"00408",
14449=>x"00408",
14450=>x"00408",
14451=>x"00408",
14452=>x"00408",
14453=>x"00408",
14454=>x"00408",
14455=>x"00408",
14456=>x"00408",
14457=>x"00408",
14458=>x"00408",
14459=>x"00408",
14460=>x"00408",
14461=>x"00408",
14462=>x"00409",
14463=>x"00409",
14464=>x"00409",
14465=>x"00409",
14466=>x"00409",
14467=>x"00409",
14468=>x"00409",
14469=>x"00409",
14470=>x"00409",
14471=>x"00409",
14472=>x"00409",
14473=>x"00409",
14474=>x"00409",
14475=>x"00409",
14476=>x"0040a",
14477=>x"0040a",
14478=>x"0040a",
14479=>x"0040a",
14480=>x"0040a",
14481=>x"0040a",
14482=>x"0040a",
14483=>x"0040a",
14484=>x"0040a",
14485=>x"0040a",
14486=>x"0040a",
14487=>x"0040a",
14488=>x"0040a",
14489=>x"0040a",
14490=>x"0040b",
14491=>x"0040b",
14492=>x"0040b",
14493=>x"0040b",
14494=>x"0040b",
14495=>x"0040b",
14496=>x"0040b",
14497=>x"0040b",
14498=>x"0040b",
14499=>x"0040b",
14500=>x"0040b",
14501=>x"0040b",
14502=>x"0040b",
14503=>x"0040b",
14504=>x"0040c",
14505=>x"0040c",
14506=>x"0040c",
14507=>x"0040c",
14508=>x"0040c",
14509=>x"0040c",
14510=>x"0040c",
14511=>x"0040c",
14512=>x"0040c",
14513=>x"0040c",
14514=>x"0040c",
14515=>x"0040c",
14516=>x"0040c",
14517=>x"0040c",
14518=>x"0040d",
14519=>x"0040d",
14520=>x"0040d",
14521=>x"0040d",
14522=>x"0040d",
14523=>x"0040d",
14524=>x"0040d",
14525=>x"0040d",
14526=>x"0040d",
14527=>x"0040d",
14528=>x"0040d",
14529=>x"0040d",
14530=>x"0040d",
14531=>x"0040d",
14532=>x"0040e",
14533=>x"0040e",
14534=>x"0040e",
14535=>x"0040e",
14536=>x"0040e",
14537=>x"0040e",
14538=>x"0040e",
14539=>x"0040e",
14540=>x"0040e",
14541=>x"0040e",
14542=>x"0040e",
14543=>x"0040e",
14544=>x"0040e",
14545=>x"0040e",
14546=>x"0040f",
14547=>x"0040f",
14548=>x"0040f",
14549=>x"0040f",
14550=>x"0040f",
14551=>x"0040f",
14552=>x"0040f",
14553=>x"0040f",
14554=>x"0040f",
14555=>x"0040f",
14556=>x"0040f",
14557=>x"0040f",
14558=>x"0040f",
14559=>x"0040f",
14560=>x"00410",
14561=>x"00410",
14562=>x"00410",
14563=>x"00410",
14564=>x"00410",
14565=>x"00410",
14566=>x"00410",
14567=>x"00410",
14568=>x"00410",
14569=>x"00410",
14570=>x"00410",
14571=>x"00410",
14572=>x"00410",
14573=>x"00410",
14574=>x"00411",
14575=>x"00411",
14576=>x"00411",
14577=>x"00411",
14578=>x"00411",
14579=>x"00411",
14580=>x"00411",
14581=>x"00411",
14582=>x"00411",
14583=>x"00411",
14584=>x"00411",
14585=>x"00411",
14586=>x"00411",
14587=>x"00411",
14588=>x"00412",
14589=>x"00412",
14590=>x"00412",
14591=>x"00412",
14592=>x"00412",
14593=>x"00412",
14594=>x"00412",
14595=>x"00412",
14596=>x"00412",
14597=>x"00412",
14598=>x"00412",
14599=>x"00412",
14600=>x"00412",
14601=>x"00412",
14602=>x"00413",
14603=>x"00413",
14604=>x"00413",
14605=>x"00413",
14606=>x"00413",
14607=>x"00413",
14608=>x"00413",
14609=>x"00413",
14610=>x"00413",
14611=>x"00413",
14612=>x"00413",
14613=>x"00413",
14614=>x"00413",
14615=>x"00413",
14616=>x"00414",
14617=>x"00414",
14618=>x"00414",
14619=>x"00414",
14620=>x"00414",
14621=>x"00414",
14622=>x"00414",
14623=>x"00414",
14624=>x"00414",
14625=>x"00414",
14626=>x"00414",
14627=>x"00414",
14628=>x"00414",
14629=>x"00414",
14630=>x"00415",
14631=>x"00415",
14632=>x"00415",
14633=>x"00415",
14634=>x"00415",
14635=>x"00415",
14636=>x"00415",
14637=>x"00415",
14638=>x"00415",
14639=>x"00415",
14640=>x"00415",
14641=>x"00415",
14642=>x"00415",
14643=>x"00415",
14644=>x"00416",
14645=>x"00416",
14646=>x"00416",
14647=>x"00416",
14648=>x"00416",
14649=>x"00416",
14650=>x"00416",
14651=>x"00416",
14652=>x"00416",
14653=>x"00416",
14654=>x"00416",
14655=>x"00416",
14656=>x"00416",
14657=>x"00416",
14658=>x"00417",
14659=>x"00417",
14660=>x"00417",
14661=>x"00417",
14662=>x"00417",
14663=>x"00417",
14664=>x"00417",
14665=>x"00417",
14666=>x"00417",
14667=>x"00417",
14668=>x"00417",
14669=>x"00417",
14670=>x"00417",
14671=>x"00417",
14672=>x"00418",
14673=>x"00418",
14674=>x"00418",
14675=>x"00418",
14676=>x"00418",
14677=>x"00418",
14678=>x"00418",
14679=>x"00418",
14680=>x"00418",
14681=>x"00418",
14682=>x"00418",
14683=>x"00418",
14684=>x"00418",
14685=>x"00418",
14686=>x"00419",
14687=>x"00419",
14688=>x"00419",
14689=>x"00419",
14690=>x"00419",
14691=>x"00419",
14692=>x"00419",
14693=>x"00419",
14694=>x"00419",
14695=>x"00419",
14696=>x"00419",
14697=>x"00419",
14698=>x"00419",
14699=>x"00419",
14700=>x"0041a",
14701=>x"0041a",
14702=>x"0041a",
14703=>x"0041a",
14704=>x"0041a",
14705=>x"0041a",
14706=>x"0041a",
14707=>x"0041a",
14708=>x"0041a",
14709=>x"0041a",
14710=>x"0041a",
14711=>x"0041a",
14712=>x"0041a",
14713=>x"0041a",
14714=>x"0041b",
14715=>x"0041b",
14716=>x"0041b",
14717=>x"0041b",
14718=>x"0041b",
14719=>x"0041b",
14720=>x"0041b",
14721=>x"0041b",
14722=>x"0041b",
14723=>x"0041b",
14724=>x"0041b",
14725=>x"0041b",
14726=>x"0041b",
14727=>x"0041b",
14728=>x"0041c",
14729=>x"0041c",
14730=>x"0041c",
14731=>x"0041c",
14732=>x"0041c",
14733=>x"0041c",
14734=>x"0041c",
14735=>x"0041c",
14736=>x"0041c",
14737=>x"0041c",
14738=>x"0041c",
14739=>x"0041c",
14740=>x"0041c",
14741=>x"0041c",
14742=>x"0041d",
14743=>x"0041d",
14744=>x"0041d",
14745=>x"0041d",
14746=>x"0041d",
14747=>x"0041d",
14748=>x"0041d",
14749=>x"0041d",
14750=>x"0041d",
14751=>x"0041d",
14752=>x"0041d",
14753=>x"0041d",
14754=>x"0041d",
14755=>x"0041d",
14756=>x"0041e",
14757=>x"0041e",
14758=>x"0041e",
14759=>x"0041e",
14760=>x"0041e",
14761=>x"0041e",
14762=>x"0041e",
14763=>x"0041e",
14764=>x"0041e",
14765=>x"0041e",
14766=>x"0041e",
14767=>x"0041e",
14768=>x"0041e",
14769=>x"0041e",
14770=>x"0041f",
14771=>x"0041f",
14772=>x"0041f",
14773=>x"0041f",
14774=>x"0041f",
14775=>x"0041f",
14776=>x"0041f",
14777=>x"0041f",
14778=>x"0041f",
14779=>x"0041f",
14780=>x"0041f",
14781=>x"0041f",
14782=>x"0041f",
14783=>x"0041f",
14784=>x"00420",
14785=>x"00420",
14786=>x"00420",
14787=>x"00420",
14788=>x"00420",
14789=>x"00420",
14790=>x"00420",
14791=>x"00420",
14792=>x"00420",
14793=>x"00420",
14794=>x"00420",
14795=>x"00420",
14796=>x"00420",
14797=>x"00420",
14798=>x"00421",
14799=>x"00421",
14800=>x"00421",
14801=>x"00421",
14802=>x"00421",
14803=>x"00421",
14804=>x"00421",
14805=>x"00421",
14806=>x"00421",
14807=>x"00421",
14808=>x"00421",
14809=>x"00421",
14810=>x"00421",
14811=>x"00421",
14812=>x"00422",
14813=>x"00422",
14814=>x"00422",
14815=>x"00422",
14816=>x"00422",
14817=>x"00422",
14818=>x"00422",
14819=>x"00422",
14820=>x"00422",
14821=>x"00422",
14822=>x"00422",
14823=>x"00422",
14824=>x"00422",
14825=>x"00422",
14826=>x"00423",
14827=>x"00423",
14828=>x"00423",
14829=>x"00423",
14830=>x"00423",
14831=>x"00423",
14832=>x"00423",
14833=>x"00423",
14834=>x"00423",
14835=>x"00423",
14836=>x"00423",
14837=>x"00423",
14838=>x"00423",
14839=>x"00423",
14840=>x"00424",
14841=>x"00424",
14842=>x"00424",
14843=>x"00424",
14844=>x"00424",
14845=>x"00424",
14846=>x"00424",
14847=>x"00424",
14848=>x"00424",
14849=>x"00424",
14850=>x"00424",
14851=>x"00424",
14852=>x"00424",
14853=>x"00424",
14854=>x"00425",
14855=>x"00425",
14856=>x"00425",
14857=>x"00425",
14858=>x"00425",
14859=>x"00425",
14860=>x"00425",
14861=>x"00425",
14862=>x"00425",
14863=>x"00425",
14864=>x"00425",
14865=>x"00425",
14866=>x"00425",
14867=>x"00425",
14868=>x"00426",
14869=>x"00426",
14870=>x"00426",
14871=>x"00426",
14872=>x"00426",
14873=>x"00426",
14874=>x"00426",
14875=>x"00426",
14876=>x"00426",
14877=>x"00426",
14878=>x"00426",
14879=>x"00426",
14880=>x"00426",
14881=>x"00426",
14882=>x"00427",
14883=>x"00427",
14884=>x"00427",
14885=>x"00427",
14886=>x"00427",
14887=>x"00427",
14888=>x"00427",
14889=>x"00427",
14890=>x"00427",
14891=>x"00427",
14892=>x"00427",
14893=>x"00427",
14894=>x"00427",
14895=>x"00427",
14896=>x"00428",
14897=>x"00428",
14898=>x"00428",
14899=>x"00428",
14900=>x"00428",
14901=>x"00428",
14902=>x"00428",
14903=>x"00428",
14904=>x"00428",
14905=>x"00428",
14906=>x"00428",
14907=>x"00428",
14908=>x"00428",
14909=>x"00428",
14910=>x"00429",
14911=>x"00429",
14912=>x"00429",
14913=>x"00429",
14914=>x"00429",
14915=>x"00429",
14916=>x"00429",
14917=>x"00429",
14918=>x"00429",
14919=>x"00429",
14920=>x"00429",
14921=>x"00429",
14922=>x"00429",
14923=>x"00429",
14924=>x"0042a",
14925=>x"0042a",
14926=>x"0042a",
14927=>x"0042a",
14928=>x"0042a",
14929=>x"0042a",
14930=>x"0042a",
14931=>x"0042a",
14932=>x"0042a",
14933=>x"0042a",
14934=>x"0042a",
14935=>x"0042a",
14936=>x"0042a",
14937=>x"0042a",
14938=>x"0042b",
14939=>x"0042b",
14940=>x"0042b",
14941=>x"0042b",
14942=>x"0042b",
14943=>x"0042b",
14944=>x"0042b",
14945=>x"0042b",
14946=>x"0042b",
14947=>x"0042b",
14948=>x"0042b",
14949=>x"0042b",
14950=>x"0042b",
14951=>x"0042b",
14952=>x"0042c",
14953=>x"0042c",
14954=>x"0042c",
14955=>x"0042c",
14956=>x"0042c",
14957=>x"0042c",
14958=>x"0042c",
14959=>x"0042c",
14960=>x"0042c",
14961=>x"0042c",
14962=>x"0042c",
14963=>x"0042c",
14964=>x"0042c",
14965=>x"0042c",
14966=>x"0042d",
14967=>x"0042d",
14968=>x"0042d",
14969=>x"0042d",
14970=>x"0042d",
14971=>x"0042d",
14972=>x"0042d",
14973=>x"0042d",
14974=>x"0042d",
14975=>x"0042d",
14976=>x"0042d",
14977=>x"0042d",
14978=>x"0042d",
14979=>x"0042d",
14980=>x"0042e",
14981=>x"0042e",
14982=>x"0042e",
14983=>x"0042e",
14984=>x"0042e",
14985=>x"0042e",
14986=>x"0042e",
14987=>x"0042e",
14988=>x"0042e",
14989=>x"0042e",
14990=>x"0042e",
14991=>x"0042e",
14992=>x"0042e",
14993=>x"0042e",
14994=>x"0042f",
14995=>x"0042f",
14996=>x"0042f",
14997=>x"0042f",
14998=>x"0042f",
14999=>x"0042f",

others=>x"00000"
);
begin
Cout<=memory(to_integer(unsigned(addr)));

end Behavioral;