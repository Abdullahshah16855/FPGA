library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.ALL;

entity RSI_ROM is
    Port ( addr : in STD_LOGIC_VECTOR (11 downto 0);
           Cout : out STD_LOGIC_VECTOR (19 downto 0));
end RSI_ROM;

architecture Behavioral of RSI_ROM is
type vector is Array(0 to 4095) of Std_logic_vector(19 downto 0);
Constant memory: vector:=
(
0=>x"00000",
1=>x"00000",
2=>x"00001",
3=>x"00002",
4=>x"00003",
5=>x"00003",
6=>x"00004",
7=>x"00005",
8=>x"00005",
9=>x"00006",
10=>x"00007",
11=>x"00007",
12=>x"00008",
13=>x"00009",
14=>x"00009",
15=>x"0000a",
16=>x"0000b",
17=>x"0000b",
18=>x"0000c",
19=>x"0000c",
20=>x"0000d",
21=>x"0000e",
22=>x"0000e",
23=>x"0000f",
24=>x"0000f",
25=>x"00010",
26=>x"00010",
27=>x"00011",
28=>x"00011",
29=>x"00012",
30=>x"00012",
31=>x"00013",
32=>x"00014",
33=>x"00014",
34=>x"00014",
35=>x"00015",
36=>x"00015",
37=>x"00016",
38=>x"00016",
39=>x"00017",
40=>x"00017",
41=>x"00018",
42=>x"00018",
43=>x"00019",
44=>x"00019",
45=>x"0001a",
46=>x"0001a",
47=>x"0001a",
48=>x"0001b",
49=>x"0001b",
50=>x"0001c",
51=>x"0001c",
52=>x"0001c",
53=>x"0001d",
54=>x"0001d",
55=>x"0001e",
56=>x"0001e",
57=>x"0001e",
58=>x"0001f",
59=>x"0001f",
60=>x"0001f",
61=>x"00020",
62=>x"00020",
63=>x"00020",
64=>x"00021",
65=>x"00021",
66=>x"00022",
67=>x"00022",
68=>x"00022",
69=>x"00023",
70=>x"00023",
71=>x"00023",
72=>x"00024",
73=>x"00024",
74=>x"00024",
75=>x"00024",
76=>x"00025",
77=>x"00025",
78=>x"00025",
79=>x"00026",
80=>x"00026",
81=>x"00026",
82=>x"00027",
83=>x"00027",
84=>x"00027",
85=>x"00027",
86=>x"00028",
87=>x"00028",
88=>x"00028",
89=>x"00029",
90=>x"00029",
91=>x"00029",
92=>x"00029",
93=>x"0002a",
94=>x"0002a",
95=>x"0002a",
96=>x"0002a",
97=>x"0002b",
98=>x"0002b",
99=>x"0002b",
100=>x"0002b",
101=>x"0002c",
102=>x"0002c",
103=>x"0002c",
104=>x"0002c",
105=>x"0002d",
106=>x"0002d",
107=>x"0002d",
108=>x"0002d",
109=>x"0002d",
110=>x"0002e",
111=>x"0002e",
112=>x"0002e",
113=>x"0002e",
114=>x"0002f",
115=>x"0002f",
116=>x"0002f",
117=>x"0002f",
118=>x"0002f",
119=>x"00030",
120=>x"00030",
121=>x"00030",
122=>x"00030",
123=>x"00031",
124=>x"00031",
125=>x"00031",
126=>x"00031",
127=>x"00031",
128=>x"00032",
129=>x"00032",
130=>x"00032",
131=>x"00032",
132=>x"00032",
133=>x"00032",
134=>x"00033",
135=>x"00033",
136=>x"00033",
137=>x"00033",
138=>x"00033",
139=>x"00034",
140=>x"00034",
141=>x"00034",
142=>x"00034",
143=>x"00034",
144=>x"00034",
145=>x"00035",
146=>x"00035",
147=>x"00035",
148=>x"00035",
149=>x"00035",
150=>x"00035",
151=>x"00036",
152=>x"00036",
153=>x"00036",
154=>x"00036",
155=>x"00036",
156=>x"00036",
157=>x"00037",
158=>x"00037",
159=>x"00037",
160=>x"00037",
161=>x"00037",
162=>x"00037",
163=>x"00038",
164=>x"00038",
165=>x"00038",
166=>x"00038",
167=>x"00038",
168=>x"00038",
169=>x"00038",
170=>x"00039",
171=>x"00039",
172=>x"00039",
173=>x"00039",
174=>x"00039",
175=>x"00039",
176=>x"00039",
177=>x"0003a",
178=>x"0003a",
179=>x"0003a",
180=>x"0003a",
181=>x"0003a",
182=>x"0003a",
183=>x"0003a",
184=>x"0003a",
185=>x"0003b",
186=>x"0003b",
187=>x"0003b",
188=>x"0003b",
189=>x"0003b",
190=>x"0003b",
191=>x"0003b",
192=>x"0003c",
193=>x"0003c",
194=>x"0003c",
195=>x"0003c",
196=>x"0003c",
197=>x"0003c",
198=>x"0003c",
199=>x"0003c",
200=>x"0003c",
201=>x"0003d",
202=>x"0003d",
203=>x"0003d",
204=>x"0003d",
205=>x"0003d",
206=>x"0003d",
207=>x"0003d",
208=>x"0003d",
209=>x"0003e",
210=>x"0003e",
211=>x"0003e",
212=>x"0003e",
213=>x"0003e",
214=>x"0003e",
215=>x"0003e",
216=>x"0003e",
217=>x"0003e",
218=>x"0003f",
219=>x"0003f",
220=>x"0003f",
221=>x"0003f",
222=>x"0003f",
223=>x"0003f",
224=>x"0003f",
225=>x"0003f",
226=>x"0003f",
227=>x"0003f",
228=>x"00040",
229=>x"00040",
230=>x"00040",
231=>x"00040",
232=>x"00040",
233=>x"00040",
234=>x"00040",
235=>x"00040",
236=>x"00040",
237=>x"00040",
238=>x"00041",
239=>x"00041",
240=>x"00041",
241=>x"00041",
242=>x"00041",
243=>x"00041",
244=>x"00041",
245=>x"00041",
246=>x"00041",
247=>x"00041",
248=>x"00041",
249=>x"00042",
250=>x"00042",
251=>x"00042",
252=>x"00042",
253=>x"00042",
254=>x"00042",
255=>x"00042",
256=>x"00042",
257=>x"00042",
258=>x"00042",
259=>x"00042",
260=>x"00043",
261=>x"00043",
262=>x"00043",
263=>x"00043",
264=>x"00043",
265=>x"00043",
266=>x"00043",
267=>x"00043",
268=>x"00043",
269=>x"00043",
270=>x"00043",
271=>x"00043",
272=>x"00044",
273=>x"00044",
274=>x"00044",
275=>x"00044",
276=>x"00044",
277=>x"00044",
278=>x"00044",
279=>x"00044",
280=>x"00044",
281=>x"00044",
282=>x"00044",
283=>x"00044",
284=>x"00044",
285=>x"00045",
286=>x"00045",
287=>x"00045",
288=>x"00045",
289=>x"00045",
290=>x"00045",
291=>x"00045",
292=>x"00045",
293=>x"00045",
294=>x"00045",
295=>x"00045",
296=>x"00045",
297=>x"00045",
298=>x"00045",
299=>x"00046",
300=>x"00046",
301=>x"00046",
302=>x"00046",
303=>x"00046",
304=>x"00046",
305=>x"00046",
306=>x"00046",
307=>x"00046",
308=>x"00046",
309=>x"00046",
310=>x"00046",
311=>x"00046",
312=>x"00046",
313=>x"00046",
314=>x"00047",
315=>x"00047",
316=>x"00047",
317=>x"00047",
318=>x"00047",
319=>x"00047",
320=>x"00047",
321=>x"00047",
322=>x"00047",
323=>x"00047",
324=>x"00047",
325=>x"00047",
326=>x"00047",
327=>x"00047",
328=>x"00047",
329=>x"00047",
330=>x"00048",
331=>x"00048",
332=>x"00048",
333=>x"00048",
334=>x"00048",
335=>x"00048",
336=>x"00048",
337=>x"00048",
338=>x"00048",
339=>x"00048",
340=>x"00048",
341=>x"00048",
342=>x"00048",
343=>x"00048",
344=>x"00048",
345=>x"00048",
346=>x"00048",
347=>x"00049",
348=>x"00049",
349=>x"00049",
350=>x"00049",
351=>x"00049",
352=>x"00049",
353=>x"00049",
354=>x"00049",
355=>x"00049",
356=>x"00049",
357=>x"00049",
358=>x"00049",
359=>x"00049",
360=>x"00049",
361=>x"00049",
362=>x"00049",
363=>x"00049",
364=>x"00049",
365=>x"0004a",
366=>x"0004a",
367=>x"0004a",
368=>x"0004a",
369=>x"0004a",
370=>x"0004a",
371=>x"0004a",
372=>x"0004a",
373=>x"0004a",
374=>x"0004a",
375=>x"0004a",
376=>x"0004a",
377=>x"0004a",
378=>x"0004a",
379=>x"0004a",
380=>x"0004a",
381=>x"0004a",
382=>x"0004a",
383=>x"0004a",
384=>x"0004b",
385=>x"0004b",
386=>x"0004b",
387=>x"0004b",
388=>x"0004b",
389=>x"0004b",
390=>x"0004b",
391=>x"0004b",
392=>x"0004b",
393=>x"0004b",
394=>x"0004b",
395=>x"0004b",
396=>x"0004b",
397=>x"0004b",
398=>x"0004b",
399=>x"0004b",
400=>x"0004b",
401=>x"0004b",
402=>x"0004b",
403=>x"0004b",
404=>x"0004b",
405=>x"0004b",
406=>x"0004c",
407=>x"0004c",
408=>x"0004c",
409=>x"0004c",
410=>x"0004c",
411=>x"0004c",
412=>x"0004c",
413=>x"0004c",
414=>x"0004c",
415=>x"0004c",
416=>x"0004c",
417=>x"0004c",
418=>x"0004c",
419=>x"0004c",
420=>x"0004c",
421=>x"0004c",
422=>x"0004c",
423=>x"0004c",
424=>x"0004c",
425=>x"0004c",
426=>x"0004c",
427=>x"0004c",
428=>x"0004c",
429=>x"0004d",
430=>x"0004d",
431=>x"0004d",
432=>x"0004d",
433=>x"0004d",
434=>x"0004d",
435=>x"0004d",
436=>x"0004d",
437=>x"0004d",
438=>x"0004d",
439=>x"0004d",
440=>x"0004d",
441=>x"0004d",
442=>x"0004d",
443=>x"0004d",
444=>x"0004d",
445=>x"0004d",
446=>x"0004d",
447=>x"0004d",
448=>x"0004d",
449=>x"0004d",
450=>x"0004d",
451=>x"0004d",
452=>x"0004d",
453=>x"0004d",
454=>x"0004e",
455=>x"0004e",
456=>x"0004e",
457=>x"0004e",
458=>x"0004e",
459=>x"0004e",
460=>x"0004e",
461=>x"0004e",
462=>x"0004e",
463=>x"0004e",
464=>x"0004e",
465=>x"0004e",
466=>x"0004e",
467=>x"0004e",
468=>x"0004e",
469=>x"0004e",
470=>x"0004e",
471=>x"0004e",
472=>x"0004e",
473=>x"0004e",
474=>x"0004e",
475=>x"0004e",
476=>x"0004e",
477=>x"0004e",
478=>x"0004e",
479=>x"0004e",
480=>x"0004e",
481=>x"0004e",
482=>x"0004f",
483=>x"0004f",
484=>x"0004f",
485=>x"0004f",
486=>x"0004f",
487=>x"0004f",
488=>x"0004f",
489=>x"0004f",
490=>x"0004f",
491=>x"0004f",
492=>x"0004f",
493=>x"0004f",
494=>x"0004f",
495=>x"0004f",
496=>x"0004f",
497=>x"0004f",
498=>x"0004f",
499=>x"0004f",
500=>x"0004f",
501=>x"0004f",
502=>x"0004f",
503=>x"0004f",
504=>x"0004f",
505=>x"0004f",
506=>x"0004f",
507=>x"0004f",
508=>x"0004f",
509=>x"0004f",
510=>x"0004f",
511=>x"0004f",
512=>x"00050",
513=>x"00050",
514=>x"00050",
515=>x"00050",
516=>x"00050",
517=>x"00050",
518=>x"00050",
519=>x"00050",
520=>x"00050",
521=>x"00050",
522=>x"00050",
523=>x"00050",
524=>x"00050",
525=>x"00050",
526=>x"00050",
527=>x"00050",
528=>x"00050",
529=>x"00050",
530=>x"00050",
531=>x"00050",
532=>x"00050",
533=>x"00050",
534=>x"00050",
535=>x"00050",
536=>x"00050",
537=>x"00050",
538=>x"00050",
539=>x"00050",
540=>x"00050",
541=>x"00050",
542=>x"00050",
543=>x"00050",
544=>x"00050",
545=>x"00050",
546=>x"00051",
547=>x"00051",
548=>x"00051",
549=>x"00051",
550=>x"00051",
551=>x"00051",
552=>x"00051",
553=>x"00051",
554=>x"00051",
555=>x"00051",
556=>x"00051",
557=>x"00051",
558=>x"00051",
559=>x"00051",
560=>x"00051",
561=>x"00051",
562=>x"00051",
563=>x"00051",
564=>x"00051",
565=>x"00051",
566=>x"00051",
567=>x"00051",
568=>x"00051",
569=>x"00051",
570=>x"00051",
571=>x"00051",
572=>x"00051",
573=>x"00051",
574=>x"00051",
575=>x"00051",
576=>x"00051",
577=>x"00051",
578=>x"00051",
579=>x"00051",
580=>x"00051",
581=>x"00051",
582=>x"00051",
583=>x"00051",
584=>x"00052",
585=>x"00052",
586=>x"00052",
587=>x"00052",
588=>x"00052",
589=>x"00052",
590=>x"00052",
591=>x"00052",
592=>x"00052",
593=>x"00052",
594=>x"00052",
595=>x"00052",
596=>x"00052",
597=>x"00052",
598=>x"00052",
599=>x"00052",
600=>x"00052",
601=>x"00052",
602=>x"00052",
603=>x"00052",
604=>x"00052",
605=>x"00052",
606=>x"00052",
607=>x"00052",
608=>x"00052",
609=>x"00052",
610=>x"00052",
611=>x"00052",
612=>x"00052",
613=>x"00052",
614=>x"00052",
615=>x"00052",
616=>x"00052",
617=>x"00052",
618=>x"00052",
619=>x"00052",
620=>x"00052",
621=>x"00052",
622=>x"00052",
623=>x"00052",
624=>x"00052",
625=>x"00053",
626=>x"00053",
627=>x"00053",
628=>x"00053",
629=>x"00053",
630=>x"00053",
631=>x"00053",
632=>x"00053",
633=>x"00053",
634=>x"00053",
635=>x"00053",
636=>x"00053",
637=>x"00053",
638=>x"00053",
639=>x"00053",
640=>x"00053",
641=>x"00053",
642=>x"00053",
643=>x"00053",
644=>x"00053",
645=>x"00053",
646=>x"00053",
647=>x"00053",
648=>x"00053",
649=>x"00053",
650=>x"00053",
651=>x"00053",
652=>x"00053",
653=>x"00053",
654=>x"00053",
655=>x"00053",
656=>x"00053",
657=>x"00053",
658=>x"00053",
659=>x"00053",
660=>x"00053",
661=>x"00053",
662=>x"00053",
663=>x"00053",
664=>x"00053",
665=>x"00053",
666=>x"00053",
667=>x"00053",
668=>x"00053",
669=>x"00053",
670=>x"00053",
671=>x"00053",
672=>x"00054",
673=>x"00054",
674=>x"00054",
675=>x"00054",
676=>x"00054",
677=>x"00054",
678=>x"00054",
679=>x"00054",
680=>x"00054",
681=>x"00054",
682=>x"00054",
683=>x"00054",
684=>x"00054",
685=>x"00054",
686=>x"00054",
687=>x"00054",
688=>x"00054",
689=>x"00054",
690=>x"00054",
691=>x"00054",
692=>x"00054",
693=>x"00054",
694=>x"00054",
695=>x"00054",
696=>x"00054",
697=>x"00054",
698=>x"00054",
699=>x"00054",
700=>x"00054",
701=>x"00054",
702=>x"00054",
703=>x"00054",
704=>x"00054",
705=>x"00054",
706=>x"00054",
707=>x"00054",
708=>x"00054",
709=>x"00054",
710=>x"00054",
711=>x"00054",
712=>x"00054",
713=>x"00054",
714=>x"00054",
715=>x"00054",
716=>x"00054",
717=>x"00054",
718=>x"00054",
719=>x"00054",
720=>x"00054",
721=>x"00054",
722=>x"00054",
723=>x"00054",
724=>x"00054",
725=>x"00054",
726=>x"00055",
727=>x"00055",
728=>x"00055",
729=>x"00055",
730=>x"00055",
731=>x"00055",
732=>x"00055",
733=>x"00055",
734=>x"00055",
735=>x"00055",
736=>x"00055",
737=>x"00055",
738=>x"00055",
739=>x"00055",
740=>x"00055",
741=>x"00055",
742=>x"00055",
743=>x"00055",
744=>x"00055",
745=>x"00055",
746=>x"00055",
747=>x"00055",
748=>x"00055",
749=>x"00055",
750=>x"00055",
751=>x"00055",
752=>x"00055",
753=>x"00055",
754=>x"00055",
755=>x"00055",
756=>x"00055",
757=>x"00055",
758=>x"00055",
759=>x"00055",
760=>x"00055",
761=>x"00055",
762=>x"00055",
763=>x"00055",
764=>x"00055",
765=>x"00055",
766=>x"00055",
767=>x"00055",
768=>x"00055",
769=>x"00055",
770=>x"00055",
771=>x"00055",
772=>x"00055",
773=>x"00055",
774=>x"00055",
775=>x"00055",
776=>x"00055",
777=>x"00055",
778=>x"00055",
779=>x"00055",
780=>x"00055",
781=>x"00055",
782=>x"00055",
783=>x"00055",
784=>x"00055",
785=>x"00055",
786=>x"00055",
787=>x"00056",
788=>x"00056",
789=>x"00056",
790=>x"00056",
791=>x"00056",
792=>x"00056",
793=>x"00056",
794=>x"00056",
795=>x"00056",
796=>x"00056",
797=>x"00056",
798=>x"00056",
799=>x"00056",
800=>x"00056",
801=>x"00056",
802=>x"00056",
803=>x"00056",
804=>x"00056",
805=>x"00056",
806=>x"00056",
807=>x"00056",
808=>x"00056",
809=>x"00056",
810=>x"00056",
811=>x"00056",
812=>x"00056",
813=>x"00056",
814=>x"00056",
815=>x"00056",
816=>x"00056",
817=>x"00056",
818=>x"00056",
819=>x"00056",
820=>x"00056",
821=>x"00056",
822=>x"00056",
823=>x"00056",
824=>x"00056",
825=>x"00056",
826=>x"00056",
827=>x"00056",
828=>x"00056",
829=>x"00056",
830=>x"00056",
831=>x"00056",
832=>x"00056",
833=>x"00056",
834=>x"00056",
835=>x"00056",
836=>x"00056",
837=>x"00056",
838=>x"00056",
839=>x"00056",
840=>x"00056",
841=>x"00056",
842=>x"00056",
843=>x"00056",
844=>x"00056",
845=>x"00056",
846=>x"00056",
847=>x"00056",
848=>x"00056",
849=>x"00056",
850=>x"00056",
851=>x"00056",
852=>x"00056",
853=>x"00056",
854=>x"00056",
855=>x"00056",
856=>x"00056",
857=>x"00057",
858=>x"00057",
859=>x"00057",
860=>x"00057",
861=>x"00057",
862=>x"00057",
863=>x"00057",
864=>x"00057",
865=>x"00057",
866=>x"00057",
867=>x"00057",
868=>x"00057",
869=>x"00057",
870=>x"00057",
871=>x"00057",
872=>x"00057",
873=>x"00057",
874=>x"00057",
875=>x"00057",
876=>x"00057",
877=>x"00057",
878=>x"00057",
879=>x"00057",
880=>x"00057",
881=>x"00057",
882=>x"00057",
883=>x"00057",
884=>x"00057",
885=>x"00057",
886=>x"00057",
887=>x"00057",
888=>x"00057",
889=>x"00057",
890=>x"00057",
891=>x"00057",
892=>x"00057",
893=>x"00057",
894=>x"00057",
895=>x"00057",
896=>x"00057",
897=>x"00057",
898=>x"00057",
899=>x"00057",
900=>x"00057",
901=>x"00057",
902=>x"00057",
903=>x"00057",
904=>x"00057",
905=>x"00057",
906=>x"00057",
907=>x"00057",
908=>x"00057",
909=>x"00057",
910=>x"00057",
911=>x"00057",
912=>x"00057",
913=>x"00057",
914=>x"00057",
915=>x"00057",
916=>x"00057",
917=>x"00057",
918=>x"00057",
919=>x"00057",
920=>x"00057",
921=>x"00057",
922=>x"00057",
923=>x"00057",
924=>x"00057",
925=>x"00057",
926=>x"00057",
927=>x"00057",
928=>x"00057",
929=>x"00057",
930=>x"00057",
931=>x"00057",
932=>x"00057",
933=>x"00057",
934=>x"00057",
935=>x"00057",
936=>x"00057",
937=>x"00057",
938=>x"00057",
939=>x"00058",
940=>x"00058",
941=>x"00058",
942=>x"00058",
943=>x"00058",
944=>x"00058",
945=>x"00058",
946=>x"00058",
947=>x"00058",
948=>x"00058",
949=>x"00058",
950=>x"00058",
951=>x"00058",
952=>x"00058",
953=>x"00058",
954=>x"00058",
955=>x"00058",
956=>x"00058",
957=>x"00058",
958=>x"00058",
959=>x"00058",
960=>x"00058",
961=>x"00058",
962=>x"00058",
963=>x"00058",
964=>x"00058",
965=>x"00058",
966=>x"00058",
967=>x"00058",
968=>x"00058",
969=>x"00058",
970=>x"00058",
971=>x"00058",
972=>x"00058",
973=>x"00058",
974=>x"00058",
975=>x"00058",
976=>x"00058",
977=>x"00058",
978=>x"00058",
979=>x"00058",
980=>x"00058",
981=>x"00058",
982=>x"00058",
983=>x"00058",
984=>x"00058",
985=>x"00058",
986=>x"00058",
987=>x"00058",
988=>x"00058",
989=>x"00058",
990=>x"00058",
991=>x"00058",
992=>x"00058",
993=>x"00058",
994=>x"00058",
995=>x"00058",
996=>x"00058",
997=>x"00058",
998=>x"00058",
999=>x"00058",
1000=>x"00058",
1001=>x"00058",
1002=>x"00058",
1003=>x"00058",
1004=>x"00058",
1005=>x"00058",
1006=>x"00058",
1007=>x"00058",
1008=>x"00058",
1009=>x"00058",
1010=>x"00058",
1011=>x"00058",
1012=>x"00058",
1013=>x"00058",
1014=>x"00058",
1015=>x"00058",
1016=>x"00058",
1017=>x"00058",
1018=>x"00058",
1019=>x"00058",
1020=>x"00058",
1021=>x"00058",
1022=>x"00058",
1023=>x"00058",
1024=>x"00058",
1025=>x"00058",
1026=>x"00058",
1027=>x"00058",
1028=>x"00058",
1029=>x"00058",
1030=>x"00058",
1031=>x"00058",
1032=>x"00058",
1033=>x"00058",
1034=>x"00058",
1035=>x"00058",
1036=>x"00059",
1037=>x"00059",
1038=>x"00059",
1039=>x"00059",
1040=>x"00059",
1041=>x"00059",
1042=>x"00059",
1043=>x"00059",
1044=>x"00059",
1045=>x"00059",
1046=>x"00059",
1047=>x"00059",
1048=>x"00059",
1049=>x"00059",
1050=>x"00059",
1051=>x"00059",
1052=>x"00059",
1053=>x"00059",
1054=>x"00059",
1055=>x"00059",
1056=>x"00059",
1057=>x"00059",
1058=>x"00059",
1059=>x"00059",
1060=>x"00059",
1061=>x"00059",
1062=>x"00059",
1063=>x"00059",
1064=>x"00059",
1065=>x"00059",
1066=>x"00059",
1067=>x"00059",
1068=>x"00059",
1069=>x"00059",
1070=>x"00059",
1071=>x"00059",
1072=>x"00059",
1073=>x"00059",
1074=>x"00059",
1075=>x"00059",
1076=>x"00059",
1077=>x"00059",
1078=>x"00059",
1079=>x"00059",
1080=>x"00059",
1081=>x"00059",
1082=>x"00059",
1083=>x"00059",
1084=>x"00059",
1085=>x"00059",
1086=>x"00059",
1087=>x"00059",
1088=>x"00059",
1089=>x"00059",
1090=>x"00059",
1091=>x"00059",
1092=>x"00059",
1093=>x"00059",
1094=>x"00059",
1095=>x"00059",
1096=>x"00059",
1097=>x"00059",
1098=>x"00059",
1099=>x"00059",
1100=>x"00059",
1101=>x"00059",
1102=>x"00059",
1103=>x"00059",
1104=>x"00059",
1105=>x"00059",
1106=>x"00059",
1107=>x"00059",
1108=>x"00059",
1109=>x"00059",
1110=>x"00059",
1111=>x"00059",
1112=>x"00059",
1113=>x"00059",
1114=>x"00059",
1115=>x"00059",
1116=>x"00059",
1117=>x"00059",
1118=>x"00059",
1119=>x"00059",
1120=>x"00059",
1121=>x"00059",
1122=>x"00059",
1123=>x"00059",
1124=>x"00059",
1125=>x"00059",
1126=>x"00059",
1127=>x"00059",
1128=>x"00059",
1129=>x"00059",
1130=>x"00059",
1131=>x"00059",
1132=>x"00059",
1133=>x"00059",
1134=>x"00059",
1135=>x"00059",
1136=>x"00059",
1137=>x"00059",
1138=>x"00059",
1139=>x"00059",
1140=>x"00059",
1141=>x"00059",
1142=>x"00059",
1143=>x"00059",
1144=>x"00059",
1145=>x"00059",
1146=>x"00059",
1147=>x"00059",
1148=>x"00059",
1149=>x"00059",
1150=>x"00059",
1151=>x"00059",
1152=>x"0005a",
1153=>x"0005a",
1154=>x"0005a",
1155=>x"0005a",
1156=>x"0005a",
1157=>x"0005a",
1158=>x"0005a",
1159=>x"0005a",
1160=>x"0005a",
1161=>x"0005a",
1162=>x"0005a",
1163=>x"0005a",
1164=>x"0005a",
1165=>x"0005a",
1166=>x"0005a",
1167=>x"0005a",
1168=>x"0005a",
1169=>x"0005a",
1170=>x"0005a",
1171=>x"0005a",
1172=>x"0005a",
1173=>x"0005a",
1174=>x"0005a",
1175=>x"0005a",
1176=>x"0005a",
1177=>x"0005a",
1178=>x"0005a",
1179=>x"0005a",
1180=>x"0005a",
1181=>x"0005a",
1182=>x"0005a",
1183=>x"0005a",
1184=>x"0005a",
1185=>x"0005a",
1186=>x"0005a",
1187=>x"0005a",
1188=>x"0005a",
1189=>x"0005a",
1190=>x"0005a",
1191=>x"0005a",
1192=>x"0005a",
1193=>x"0005a",
1194=>x"0005a",
1195=>x"0005a",
1196=>x"0005a",
1197=>x"0005a",
1198=>x"0005a",
1199=>x"0005a",
1200=>x"0005a",
1201=>x"0005a",
1202=>x"0005a",
1203=>x"0005a",
1204=>x"0005a",
1205=>x"0005a",
1206=>x"0005a",
1207=>x"0005a",
1208=>x"0005a",
1209=>x"0005a",
1210=>x"0005a",
1211=>x"0005a",
1212=>x"0005a",
1213=>x"0005a",
1214=>x"0005a",
1215=>x"0005a",
1216=>x"0005a",
1217=>x"0005a",
1218=>x"0005a",
1219=>x"0005a",
1220=>x"0005a",
1221=>x"0005a",
1222=>x"0005a",
1223=>x"0005a",
1224=>x"0005a",
1225=>x"0005a",
1226=>x"0005a",
1227=>x"0005a",
1228=>x"0005a",
1229=>x"0005a",
1230=>x"0005a",
1231=>x"0005a",
1232=>x"0005a",
1233=>x"0005a",
1234=>x"0005a",
1235=>x"0005a",
1236=>x"0005a",
1237=>x"0005a",
1238=>x"0005a",
1239=>x"0005a",
1240=>x"0005a",
1241=>x"0005a",
1242=>x"0005a",
1243=>x"0005a",
1244=>x"0005a",
1245=>x"0005a",
1246=>x"0005a",
1247=>x"0005a",
1248=>x"0005a",
1249=>x"0005a",
1250=>x"0005a",
1251=>x"0005a",
1252=>x"0005a",
1253=>x"0005a",
1254=>x"0005a",
1255=>x"0005a",
1256=>x"0005a",
1257=>x"0005a",
1258=>x"0005a",
1259=>x"0005a",
1260=>x"0005a",
1261=>x"0005a",
1262=>x"0005a",
1263=>x"0005a",
1264=>x"0005a",
1265=>x"0005a",
1266=>x"0005a",
1267=>x"0005a",
1268=>x"0005a",
1269=>x"0005a",
1270=>x"0005a",
1271=>x"0005a",
1272=>x"0005a",
1273=>x"0005a",
1274=>x"0005a",
1275=>x"0005a",
1276=>x"0005a",
1277=>x"0005a",
1278=>x"0005a",
1279=>x"0005a",
1280=>x"0005a",
1281=>x"0005a",
1282=>x"0005a",
1283=>x"0005a",
1284=>x"0005a",
1285=>x"0005a",
1286=>x"0005a",
1287=>x"0005a",
1288=>x"0005a",
1289=>x"0005a",
1290=>x"0005a",
1291=>x"0005a",
1292=>x"0005a",
1293=>x"0005a",
1294=>x"0005a",
1295=>x"0005b",
1296=>x"0005b",
1297=>x"0005b",
1298=>x"0005b",
1299=>x"0005b",
1300=>x"0005b",
1301=>x"0005b",
1302=>x"0005b",
1303=>x"0005b",
1304=>x"0005b",
1305=>x"0005b",
1306=>x"0005b",
1307=>x"0005b",
1308=>x"0005b",
1309=>x"0005b",
1310=>x"0005b",
1311=>x"0005b",
1312=>x"0005b",
1313=>x"0005b",
1314=>x"0005b",
1315=>x"0005b",
1316=>x"0005b",
1317=>x"0005b",
1318=>x"0005b",
1319=>x"0005b",
1320=>x"0005b",
1321=>x"0005b",
1322=>x"0005b",
1323=>x"0005b",
1324=>x"0005b",
1325=>x"0005b",
1326=>x"0005b",
1327=>x"0005b",
1328=>x"0005b",
1329=>x"0005b",
1330=>x"0005b",
1331=>x"0005b",
1332=>x"0005b",
1333=>x"0005b",
1334=>x"0005b",
1335=>x"0005b",
1336=>x"0005b",
1337=>x"0005b",
1338=>x"0005b",
1339=>x"0005b",
1340=>x"0005b",
1341=>x"0005b",
1342=>x"0005b",
1343=>x"0005b",
1344=>x"0005b",
1345=>x"0005b",
1346=>x"0005b",
1347=>x"0005b",
1348=>x"0005b",
1349=>x"0005b",
1350=>x"0005b",
1351=>x"0005b",
1352=>x"0005b",
1353=>x"0005b",
1354=>x"0005b",
1355=>x"0005b",
1356=>x"0005b",
1357=>x"0005b",
1358=>x"0005b",
1359=>x"0005b",
1360=>x"0005b",
1361=>x"0005b",
1362=>x"0005b",
1363=>x"0005b",
1364=>x"0005b",
1365=>x"0005b",
1366=>x"0005b",
1367=>x"0005b",
1368=>x"0005b",
1369=>x"0005b",
1370=>x"0005b",
1371=>x"0005b",
1372=>x"0005b",
1373=>x"0005b",
1374=>x"0005b",
1375=>x"0005b",
1376=>x"0005b",
1377=>x"0005b",
1378=>x"0005b",
1379=>x"0005b",
1380=>x"0005b",
1381=>x"0005b",
1382=>x"0005b",
1383=>x"0005b",
1384=>x"0005b",
1385=>x"0005b",
1386=>x"0005b",
1387=>x"0005b",
1388=>x"0005b",
1389=>x"0005b",
1390=>x"0005b",
1391=>x"0005b",
1392=>x"0005b",
1393=>x"0005b",
1394=>x"0005b",
1395=>x"0005b",
1396=>x"0005b",
1397=>x"0005b",
1398=>x"0005b",
1399=>x"0005b",
1400=>x"0005b",
1401=>x"0005b",
1402=>x"0005b",
1403=>x"0005b",
1404=>x"0005b",
1405=>x"0005b",
1406=>x"0005b",
1407=>x"0005b",
1408=>x"0005b",
1409=>x"0005b",
1410=>x"0005b",
1411=>x"0005b",
1412=>x"0005b",
1413=>x"0005b",
1414=>x"0005b",
1415=>x"0005b",
1416=>x"0005b",
1417=>x"0005b",
1418=>x"0005b",
1419=>x"0005b",
1420=>x"0005b",
1421=>x"0005b",
1422=>x"0005b",
1423=>x"0005b",
1424=>x"0005b",
1425=>x"0005b",
1426=>x"0005b",
1427=>x"0005b",
1428=>x"0005b",
1429=>x"0005b",
1430=>x"0005b",
1431=>x"0005b",
1432=>x"0005b",
1433=>x"0005b",
1434=>x"0005b",
1435=>x"0005b",
1436=>x"0005b",
1437=>x"0005b",
1438=>x"0005b",
1439=>x"0005b",
1440=>x"0005b",
1441=>x"0005b",
1442=>x"0005b",
1443=>x"0005b",
1444=>x"0005b",
1445=>x"0005b",
1446=>x"0005b",
1447=>x"0005b",
1448=>x"0005b",
1449=>x"0005b",
1450=>x"0005b",
1451=>x"0005b",
1452=>x"0005b",
1453=>x"0005b",
1454=>x"0005b",
1455=>x"0005b",
1456=>x"0005b",
1457=>x"0005b",
1458=>x"0005b",
1459=>x"0005b",
1460=>x"0005b",
1461=>x"0005b",
1462=>x"0005b",
1463=>x"0005b",
1464=>x"0005b",
1465=>x"0005b",
1466=>x"0005b",
1467=>x"0005b",
1468=>x"0005b",
1469=>x"0005b",
1470=>x"0005b",
1471=>x"0005b",
1472=>x"0005c",
1473=>x"0005c",
1474=>x"0005c",
1475=>x"0005c",
1476=>x"0005c",
1477=>x"0005c",
1478=>x"0005c",
1479=>x"0005c",
1480=>x"0005c",
1481=>x"0005c",
1482=>x"0005c",
1483=>x"0005c",
1484=>x"0005c",
1485=>x"0005c",
1486=>x"0005c",
1487=>x"0005c",
1488=>x"0005c",
1489=>x"0005c",
1490=>x"0005c",
1491=>x"0005c",
1492=>x"0005c",
1493=>x"0005c",
1494=>x"0005c",
1495=>x"0005c",
1496=>x"0005c",
1497=>x"0005c",
1498=>x"0005c",
1499=>x"0005c",
1500=>x"0005c",
1501=>x"0005c",
1502=>x"0005c",
1503=>x"0005c",
1504=>x"0005c",
1505=>x"0005c",
1506=>x"0005c",
1507=>x"0005c",
1508=>x"0005c",
1509=>x"0005c",
1510=>x"0005c",
1511=>x"0005c",
1512=>x"0005c",
1513=>x"0005c",
1514=>x"0005c",
1515=>x"0005c",
1516=>x"0005c",
1517=>x"0005c",
1518=>x"0005c",
1519=>x"0005c",
1520=>x"0005c",
1521=>x"0005c",
1522=>x"0005c",
1523=>x"0005c",
1524=>x"0005c",
1525=>x"0005c",
1526=>x"0005c",
1527=>x"0005c",
1528=>x"0005c",
1529=>x"0005c",
1530=>x"0005c",
1531=>x"0005c",
1532=>x"0005c",
1533=>x"0005c",
1534=>x"0005c",
1535=>x"0005c",
1536=>x"0005c",
1537=>x"0005c",
1538=>x"0005c",
1539=>x"0005c",
1540=>x"0005c",
1541=>x"0005c",
1542=>x"0005c",
1543=>x"0005c",
1544=>x"0005c",
1545=>x"0005c",
1546=>x"0005c",
1547=>x"0005c",
1548=>x"0005c",
1549=>x"0005c",
1550=>x"0005c",
1551=>x"0005c",
1552=>x"0005c",
1553=>x"0005c",
1554=>x"0005c",
1555=>x"0005c",
1556=>x"0005c",
1557=>x"0005c",
1558=>x"0005c",
1559=>x"0005c",
1560=>x"0005c",
1561=>x"0005c",
1562=>x"0005c",
1563=>x"0005c",
1564=>x"0005c",
1565=>x"0005c",
1566=>x"0005c",
1567=>x"0005c",
1568=>x"0005c",
1569=>x"0005c",
1570=>x"0005c",
1571=>x"0005c",
1572=>x"0005c",
1573=>x"0005c",
1574=>x"0005c",
1575=>x"0005c",
1576=>x"0005c",
1577=>x"0005c",
1578=>x"0005c",
1579=>x"0005c",
1580=>x"0005c",
1581=>x"0005c",
1582=>x"0005c",
1583=>x"0005c",
1584=>x"0005c",
1585=>x"0005c",
1586=>x"0005c",
1587=>x"0005c",
1588=>x"0005c",
1589=>x"0005c",
1590=>x"0005c",
1591=>x"0005c",
1592=>x"0005c",
1593=>x"0005c",
1594=>x"0005c",
1595=>x"0005c",
1596=>x"0005c",
1597=>x"0005c",
1598=>x"0005c",
1599=>x"0005c",
1600=>x"0005c",
1601=>x"0005c",
1602=>x"0005c",
1603=>x"0005c",
1604=>x"0005c",
1605=>x"0005c",
1606=>x"0005c",
1607=>x"0005c",
1608=>x"0005c",
1609=>x"0005c",
1610=>x"0005c",
1611=>x"0005c",
1612=>x"0005c",
1613=>x"0005c",
1614=>x"0005c",
1615=>x"0005c",
1616=>x"0005c",
1617=>x"0005c",
1618=>x"0005c",
1619=>x"0005c",
1620=>x"0005c",
1621=>x"0005c",
1622=>x"0005c",
1623=>x"0005c",
1624=>x"0005c",
1625=>x"0005c",
1626=>x"0005c",
1627=>x"0005c",
1628=>x"0005c",
1629=>x"0005c",
1630=>x"0005c",
1631=>x"0005c",
1632=>x"0005c",
1633=>x"0005c",
1634=>x"0005c",
1635=>x"0005c",
1636=>x"0005c",
1637=>x"0005c",
1638=>x"0005c",
1639=>x"0005c",
1640=>x"0005c",
1641=>x"0005c",
1642=>x"0005c",
1643=>x"0005c",
1644=>x"0005c",
1645=>x"0005c",
1646=>x"0005c",
1647=>x"0005c",
1648=>x"0005c",
1649=>x"0005c",
1650=>x"0005c",
1651=>x"0005c",
1652=>x"0005c",
1653=>x"0005c",
1654=>x"0005c",
1655=>x"0005c",
1656=>x"0005c",
1657=>x"0005c",
1658=>x"0005c",
1659=>x"0005c",
1660=>x"0005c",
1661=>x"0005c",
1662=>x"0005c",
1663=>x"0005c",
1664=>x"0005c",
1665=>x"0005c",
1666=>x"0005c",
1667=>x"0005c",
1668=>x"0005c",
1669=>x"0005c",
1670=>x"0005c",
1671=>x"0005c",
1672=>x"0005c",
1673=>x"0005c",
1674=>x"0005c",
1675=>x"0005c",
1676=>x"0005c",
1677=>x"0005c",
1678=>x"0005c",
1679=>x"0005c",
1680=>x"0005c",
1681=>x"0005c",
1682=>x"0005c",
1683=>x"0005c",
1684=>x"0005c",
1685=>x"0005c",
1686=>x"0005c",
1687=>x"0005c",
1688=>x"0005c",
1689=>x"0005c",
1690=>x"0005c",
1691=>x"0005c",
1692=>x"0005c",
1693=>x"0005c",
1694=>x"0005c",
1695=>x"0005c",
1696=>x"0005c",
1697=>x"0005c",
1698=>x"0005c",
1699=>x"0005c",
1700=>x"0005c",
1701=>x"0005d",
1702=>x"0005d",
1703=>x"0005d",
1704=>x"0005d",
1705=>x"0005d",
1706=>x"0005d",
1707=>x"0005d",
1708=>x"0005d",
1709=>x"0005d",
1710=>x"0005d",
1711=>x"0005d",
1712=>x"0005d",
1713=>x"0005d",
1714=>x"0005d",
1715=>x"0005d",
1716=>x"0005d",
1717=>x"0005d",
1718=>x"0005d",
1719=>x"0005d",
1720=>x"0005d",
1721=>x"0005d",
1722=>x"0005d",
1723=>x"0005d",
1724=>x"0005d",
1725=>x"0005d",
1726=>x"0005d",
1727=>x"0005d",
1728=>x"0005d",
1729=>x"0005d",
1730=>x"0005d",
1731=>x"0005d",
1732=>x"0005d",
1733=>x"0005d",
1734=>x"0005d",
1735=>x"0005d",
1736=>x"0005d",
1737=>x"0005d",
1738=>x"0005d",
1739=>x"0005d",
1740=>x"0005d",
1741=>x"0005d",
1742=>x"0005d",
1743=>x"0005d",
1744=>x"0005d",
1745=>x"0005d",
1746=>x"0005d",
1747=>x"0005d",
1748=>x"0005d",
1749=>x"0005d",
1750=>x"0005d",
1751=>x"0005d",
1752=>x"0005d",
1753=>x"0005d",
1754=>x"0005d",
1755=>x"0005d",
1756=>x"0005d",
1757=>x"0005d",
1758=>x"0005d",
1759=>x"0005d",
1760=>x"0005d",
1761=>x"0005d",
1762=>x"0005d",
1763=>x"0005d",
1764=>x"0005d",
1765=>x"0005d",
1766=>x"0005d",
1767=>x"0005d",
1768=>x"0005d",
1769=>x"0005d",
1770=>x"0005d",
1771=>x"0005d",
1772=>x"0005d",
1773=>x"0005d",
1774=>x"0005d",
1775=>x"0005d",
1776=>x"0005d",
1777=>x"0005d",
1778=>x"0005d",
1779=>x"0005d",
1780=>x"0005d",
1781=>x"0005d",
1782=>x"0005d",
1783=>x"0005d",
1784=>x"0005d",
1785=>x"0005d",
1786=>x"0005d",
1787=>x"0005d",
1788=>x"0005d",
1789=>x"0005d",
1790=>x"0005d",
1791=>x"0005d",
1792=>x"0005d",
1793=>x"0005d",
1794=>x"0005d",
1795=>x"0005d",
1796=>x"0005d",
1797=>x"0005d",
1798=>x"0005d",
1799=>x"0005d",
1800=>x"0005d",
1801=>x"0005d",
1802=>x"0005d",
1803=>x"0005d",
1804=>x"0005d",
1805=>x"0005d",
1806=>x"0005d",
1807=>x"0005d",
1808=>x"0005d",
1809=>x"0005d",
1810=>x"0005d",
1811=>x"0005d",
1812=>x"0005d",
1813=>x"0005d",
1814=>x"0005d",
1815=>x"0005d",
1816=>x"0005d",
1817=>x"0005d",
1818=>x"0005d",
1819=>x"0005d",
1820=>x"0005d",
1821=>x"0005d",
1822=>x"0005d",
1823=>x"0005d",
1824=>x"0005d",
1825=>x"0005d",
1826=>x"0005d",
1827=>x"0005d",
1828=>x"0005d",
1829=>x"0005d",
1830=>x"0005d",
1831=>x"0005d",
1832=>x"0005d",
1833=>x"0005d",
1834=>x"0005d",
1835=>x"0005d",
1836=>x"0005d",
1837=>x"0005d",
1838=>x"0005d",
1839=>x"0005d",
1840=>x"0005d",
1841=>x"0005d",
1842=>x"0005d",
1843=>x"0005d",
1844=>x"0005d",
1845=>x"0005d",
1846=>x"0005d",
1847=>x"0005d",
1848=>x"0005d",
1849=>x"0005d",
1850=>x"0005d",
1851=>x"0005d",
1852=>x"0005d",
1853=>x"0005d",
1854=>x"0005d",
1855=>x"0005d",
1856=>x"0005d",
1857=>x"0005d",
1858=>x"0005d",
1859=>x"0005d",
1860=>x"0005d",
1861=>x"0005d",
1862=>x"0005d",
1863=>x"0005d",
1864=>x"0005d",
1865=>x"0005d",
1866=>x"0005d",
1867=>x"0005d",
1868=>x"0005d",
1869=>x"0005d",
1870=>x"0005d",
1871=>x"0005d",
1872=>x"0005d",
1873=>x"0005d",
1874=>x"0005d",
1875=>x"0005d",
1876=>x"0005d",
1877=>x"0005d",
1878=>x"0005d",
1879=>x"0005d",
1880=>x"0005d",
1881=>x"0005d",
1882=>x"0005d",
1883=>x"0005d",
1884=>x"0005d",
1885=>x"0005d",
1886=>x"0005d",
1887=>x"0005d",
1888=>x"0005d",
1889=>x"0005d",
1890=>x"0005d",
1891=>x"0005d",
1892=>x"0005d",
1893=>x"0005d",
1894=>x"0005d",
1895=>x"0005d",
1896=>x"0005d",
1897=>x"0005d",
1898=>x"0005d",
1899=>x"0005d",
1900=>x"0005d",
1901=>x"0005d",
1902=>x"0005d",
1903=>x"0005d",
1904=>x"0005d",
1905=>x"0005d",
1906=>x"0005d",
1907=>x"0005d",
1908=>x"0005d",
1909=>x"0005d",
1910=>x"0005d",
1911=>x"0005d",
1912=>x"0005d",
1913=>x"0005d",
1914=>x"0005d",
1915=>x"0005d",
1916=>x"0005d",
1917=>x"0005d",
1918=>x"0005d",
1919=>x"0005d",
1920=>x"0005d",
1921=>x"0005d",
1922=>x"0005d",
1923=>x"0005d",
1924=>x"0005d",
1925=>x"0005d",
1926=>x"0005d",
1927=>x"0005d",
1928=>x"0005d",
1929=>x"0005d",
1930=>x"0005d",
1931=>x"0005d",
1932=>x"0005d",
1933=>x"0005d",
1934=>x"0005d",
1935=>x"0005d",
1936=>x"0005d",
1937=>x"0005d",
1938=>x"0005d",
1939=>x"0005d",
1940=>x"0005d",
1941=>x"0005d",
1942=>x"0005d",
1943=>x"0005d",
1944=>x"0005d",
1945=>x"0005d",
1946=>x"0005d",
1947=>x"0005d",
1948=>x"0005d",
1949=>x"0005d",
1950=>x"0005d",
1951=>x"0005d",
1952=>x"0005d",
1953=>x"0005d",
1954=>x"0005d",
1955=>x"0005d",
1956=>x"0005d",
1957=>x"0005d",
1958=>x"0005d",
1959=>x"0005d",
1960=>x"0005d",
1961=>x"0005d",
1962=>x"0005d",
1963=>x"0005d",
1964=>x"0005d",
1965=>x"0005d",
1966=>x"0005d",
1967=>x"0005d",
1968=>x"0005d",
1969=>x"0005d",
1970=>x"0005d",
1971=>x"0005d",
1972=>x"0005d",
1973=>x"0005d",
1974=>x"0005d",
1975=>x"0005d",
1976=>x"0005d",
1977=>x"0005d",
1978=>x"0005d",
1979=>x"0005d",
1980=>x"0005d",
1981=>x"0005d",
1982=>x"0005d",
1983=>x"0005d",
1984=>x"0005d",
1985=>x"0005d",
1986=>x"0005d",
1987=>x"0005d",
1988=>x"0005d",
1989=>x"0005d",
1990=>x"0005d",
1991=>x"0005d",
1992=>x"0005d",
1993=>x"0005d",
1994=>x"0005d",
1995=>x"0005d",
1996=>x"0005d",
1997=>x"0005d",
1998=>x"0005d",
1999=>x"0005d",
2000=>x"0005d",
2001=>x"0005d",
2002=>x"0005d",
2003=>x"0005d",
2004=>x"0005d",
2005=>x"0005d",
2006=>x"0005e",
2007=>x"0005e",
2008=>x"0005e",
2009=>x"0005e",
2010=>x"0005e",
2011=>x"0005e",
2012=>x"0005e",
2013=>x"0005e",
2014=>x"0005e",
2015=>x"0005e",
2016=>x"0005e",
2017=>x"0005e",
2018=>x"0005e",
2019=>x"0005e",
2020=>x"0005e",
2021=>x"0005e",
2022=>x"0005e",
2023=>x"0005e",
2024=>x"0005e",
2025=>x"0005e",
2026=>x"0005e",
2027=>x"0005e",
2028=>x"0005e",
2029=>x"0005e",
2030=>x"0005e",
2031=>x"0005e",
2032=>x"0005e",
2033=>x"0005e",
2034=>x"0005e",
2035=>x"0005e",
2036=>x"0005e",
2037=>x"0005e",
2038=>x"0005e",
2039=>x"0005e",
2040=>x"0005e",
2041=>x"0005e",
2042=>x"0005e",
2043=>x"0005e",
2044=>x"0005e",
2045=>x"0005e",
2046=>x"0005e",
2047=>x"0005e",
2048=>x"0005e",
2049=>x"0005e",
2050=>x"0005e",
2051=>x"0005e",
2052=>x"0005e",
2053=>x"0005e",
2054=>x"0005e",
2055=>x"0005e",
2056=>x"0005e",
2057=>x"0005e",
2058=>x"0005e",
2059=>x"0005e",
2060=>x"0005e",
2061=>x"0005e",
2062=>x"0005e",
2063=>x"0005e",
2064=>x"0005e",
2065=>x"0005e",
2066=>x"0005e",
2067=>x"0005e",
2068=>x"0005e",
2069=>x"0005e",
2070=>x"0005e",
2071=>x"0005e",
2072=>x"0005e",
2073=>x"0005e",
2074=>x"0005e",
2075=>x"0005e",
2076=>x"0005e",
2077=>x"0005e",
2078=>x"0005e",
2079=>x"0005e",
2080=>x"0005e",
2081=>x"0005e",
2082=>x"0005e",
2083=>x"0005e",
2084=>x"0005e",
2085=>x"0005e",
2086=>x"0005e",
2087=>x"0005e",
2088=>x"0005e",
2089=>x"0005e",
2090=>x"0005e",
2091=>x"0005e",
2092=>x"0005e",
2093=>x"0005e",
2094=>x"0005e",
2095=>x"0005e",
2096=>x"0005e",
2097=>x"0005e",
2098=>x"0005e",
2099=>x"0005e",
2100=>x"0005e",
2101=>x"0005e",
2102=>x"0005e",
2103=>x"0005e",
2104=>x"0005e",
2105=>x"0005e",
2106=>x"0005e",
2107=>x"0005e",
2108=>x"0005e",
2109=>x"0005e",
2110=>x"0005e",
2111=>x"0005e",
2112=>x"0005e",
2113=>x"0005e",
2114=>x"0005e",
2115=>x"0005e",
2116=>x"0005e",
2117=>x"0005e",
2118=>x"0005e",
2119=>x"0005e",
2120=>x"0005e",
2121=>x"0005e",
2122=>x"0005e",
2123=>x"0005e",
2124=>x"0005e",
2125=>x"0005e",
2126=>x"0005e",
2127=>x"0005e",
2128=>x"0005e",
2129=>x"0005e",
2130=>x"0005e",
2131=>x"0005e",
2132=>x"0005e",
2133=>x"0005e",
2134=>x"0005e",
2135=>x"0005e",
2136=>x"0005e",
2137=>x"0005e",
2138=>x"0005e",
2139=>x"0005e",
2140=>x"0005e",
2141=>x"0005e",
2142=>x"0005e",
2143=>x"0005e",
2144=>x"0005e",
2145=>x"0005e",
2146=>x"0005e",
2147=>x"0005e",
2148=>x"0005e",
2149=>x"0005e",
2150=>x"0005e",
2151=>x"0005e",
2152=>x"0005e",
2153=>x"0005e",
2154=>x"0005e",
2155=>x"0005e",
2156=>x"0005e",
2157=>x"0005e",
2158=>x"0005e",
2159=>x"0005e",
2160=>x"0005e",
2161=>x"0005e",
2162=>x"0005e",
2163=>x"0005e",
2164=>x"0005e",
2165=>x"0005e",
2166=>x"0005e",
2167=>x"0005e",
2168=>x"0005e",
2169=>x"0005e",
2170=>x"0005e",
2171=>x"0005e",
2172=>x"0005e",
2173=>x"0005e",
2174=>x"0005e",
2175=>x"0005e",
2176=>x"0005e",
2177=>x"0005e",
2178=>x"0005e",
2179=>x"0005e",
2180=>x"0005e",
2181=>x"0005e",
2182=>x"0005e",
2183=>x"0005e",
2184=>x"0005e",
2185=>x"0005e",
2186=>x"0005e",
2187=>x"0005e",
2188=>x"0005e",
2189=>x"0005e",
2190=>x"0005e",
2191=>x"0005e",
2192=>x"0005e",
2193=>x"0005e",
2194=>x"0005e",
2195=>x"0005e",
2196=>x"0005e",
2197=>x"0005e",
2198=>x"0005e",
2199=>x"0005e",
2200=>x"0005e",
2201=>x"0005e",
2202=>x"0005e",
2203=>x"0005e",
2204=>x"0005e",
2205=>x"0005e",
2206=>x"0005e",
2207=>x"0005e",
2208=>x"0005e",
2209=>x"0005e",
2210=>x"0005e",
2211=>x"0005e",
2212=>x"0005e",
2213=>x"0005e",
2214=>x"0005e",
2215=>x"0005e",
2216=>x"0005e",
2217=>x"0005e",
2218=>x"0005e",
2219=>x"0005e",
2220=>x"0005e",
2221=>x"0005e",
2222=>x"0005e",
2223=>x"0005e",
2224=>x"0005e",
2225=>x"0005e",
2226=>x"0005e",
2227=>x"0005e",
2228=>x"0005e",
2229=>x"0005e",
2230=>x"0005e",
2231=>x"0005e",
2232=>x"0005e",
2233=>x"0005e",
2234=>x"0005e",
2235=>x"0005e",
2236=>x"0005e",
2237=>x"0005e",
2238=>x"0005e",
2239=>x"0005e",
2240=>x"0005e",
2241=>x"0005e",
2242=>x"0005e",
2243=>x"0005e",
2244=>x"0005e",
2245=>x"0005e",
2246=>x"0005e",
2247=>x"0005e",
2248=>x"0005e",
2249=>x"0005e",
2250=>x"0005e",
2251=>x"0005e",
2252=>x"0005e",
2253=>x"0005e",
2254=>x"0005e",
2255=>x"0005e",
2256=>x"0005e",
2257=>x"0005e",
2258=>x"0005e",
2259=>x"0005e",
2260=>x"0005e",
2261=>x"0005e",
2262=>x"0005e",
2263=>x"0005e",
2264=>x"0005e",
2265=>x"0005e",
2266=>x"0005e",
2267=>x"0005e",
2268=>x"0005e",
2269=>x"0005e",
2270=>x"0005e",
2271=>x"0005e",
2272=>x"0005e",
2273=>x"0005e",
2274=>x"0005e",
2275=>x"0005e",
2276=>x"0005e",
2277=>x"0005e",
2278=>x"0005e",
2279=>x"0005e",
2280=>x"0005e",
2281=>x"0005e",
2282=>x"0005e",
2283=>x"0005e",
2284=>x"0005e",
2285=>x"0005e",
2286=>x"0005e",
2287=>x"0005e",
2288=>x"0005e",
2289=>x"0005e",
2290=>x"0005e",
2291=>x"0005e",
2292=>x"0005e",
2293=>x"0005e",
2294=>x"0005e",
2295=>x"0005e",
2296=>x"0005e",
2297=>x"0005e",
2298=>x"0005e",
2299=>x"0005e",
2300=>x"0005e",
2301=>x"0005e",
2302=>x"0005e",
2303=>x"0005e",
2304=>x"0005e",
2305=>x"0005e",
2306=>x"0005e",
2307=>x"0005e",
2308=>x"0005e",
2309=>x"0005e",
2310=>x"0005e",
2311=>x"0005e",
2312=>x"0005e",
2313=>x"0005e",
2314=>x"0005e",
2315=>x"0005e",
2316=>x"0005e",
2317=>x"0005e",
2318=>x"0005e",
2319=>x"0005e",
2320=>x"0005e",
2321=>x"0005e",
2322=>x"0005e",
2323=>x"0005e",
2324=>x"0005e",
2325=>x"0005e",
2326=>x"0005e",
2327=>x"0005e",
2328=>x"0005e",
2329=>x"0005e",
2330=>x"0005e",
2331=>x"0005e",
2332=>x"0005e",
2333=>x"0005e",
2334=>x"0005e",
2335=>x"0005e",
2336=>x"0005e",
2337=>x"0005e",
2338=>x"0005e",
2339=>x"0005e",
2340=>x"0005e",
2341=>x"0005e",
2342=>x"0005e",
2343=>x"0005e",
2344=>x"0005e",
2345=>x"0005e",
2346=>x"0005e",
2347=>x"0005e",
2348=>x"0005e",
2349=>x"0005e",
2350=>x"0005e",
2351=>x"0005e",
2352=>x"0005e",
2353=>x"0005e",
2354=>x"0005e",
2355=>x"0005e",
2356=>x"0005e",
2357=>x"0005e",
2358=>x"0005e",
2359=>x"0005e",
2360=>x"0005e",
2361=>x"0005e",
2362=>x"0005e",
2363=>x"0005e",
2364=>x"0005e",
2365=>x"0005e",
2366=>x"0005e",
2367=>x"0005e",
2368=>x"0005e",
2369=>x"0005e",
2370=>x"0005e",
2371=>x"0005e",
2372=>x"0005e",
2373=>x"0005e",
2374=>x"0005e",
2375=>x"0005e",
2376=>x"0005e",
2377=>x"0005e",
2378=>x"0005e",
2379=>x"0005e",
2380=>x"0005e",
2381=>x"0005e",
2382=>x"0005e",
2383=>x"0005e",
2384=>x"0005e",
2385=>x"0005e",
2386=>x"0005e",
2387=>x"0005e",
2388=>x"0005e",
2389=>x"0005e",
2390=>x"0005e",
2391=>x"0005e",
2392=>x"0005e",
2393=>x"0005e",
2394=>x"0005e",
2395=>x"0005e",
2396=>x"0005e",
2397=>x"0005e",
2398=>x"0005e",
2399=>x"0005e",
2400=>x"0005e",
2401=>x"0005e",
2402=>x"0005e",
2403=>x"0005e",
2404=>x"0005e",
2405=>x"0005e",
2406=>x"0005e",
2407=>x"0005e",
2408=>x"0005e",
2409=>x"0005e",
2410=>x"0005e",
2411=>x"0005e",
2412=>x"0005e",
2413=>x"0005e",
2414=>x"0005e",
2415=>x"0005e",
2416=>x"0005e",
2417=>x"0005e",
2418=>x"0005e",
2419=>x"0005e",
2420=>x"0005e",
2421=>x"0005e",
2422=>x"0005e",
2423=>x"0005e",
2424=>x"0005e",
2425=>x"0005e",
2426=>x"0005e",
2427=>x"0005e",
2428=>x"0005e",
2429=>x"0005e",
2430=>x"0005e",
2431=>x"0005e",
2432=>x"0005f",
2433=>x"0005f",
2434=>x"0005f",
2435=>x"0005f",
2436=>x"0005f",
2437=>x"0005f",
2438=>x"0005f",
2439=>x"0005f",
2440=>x"0005f",
2441=>x"0005f",
2442=>x"0005f",
2443=>x"0005f",
2444=>x"0005f",
2445=>x"0005f",
2446=>x"0005f",
2447=>x"0005f",
2448=>x"0005f",
2449=>x"0005f",
2450=>x"0005f",
2451=>x"0005f",
2452=>x"0005f",
2453=>x"0005f",
2454=>x"0005f",
2455=>x"0005f",
2456=>x"0005f",
2457=>x"0005f",
2458=>x"0005f",
2459=>x"0005f",
2460=>x"0005f",
2461=>x"0005f",
2462=>x"0005f",
2463=>x"0005f",
2464=>x"0005f",
2465=>x"0005f",
2466=>x"0005f",
2467=>x"0005f",
2468=>x"0005f",
2469=>x"0005f",
2470=>x"0005f",
2471=>x"0005f",
2472=>x"0005f",
2473=>x"0005f",
2474=>x"0005f",
2475=>x"0005f",
2476=>x"0005f",
2477=>x"0005f",
2478=>x"0005f",
2479=>x"0005f",
2480=>x"0005f",
2481=>x"0005f",
2482=>x"0005f",
2483=>x"0005f",
2484=>x"0005f",
2485=>x"0005f",
2486=>x"0005f",
2487=>x"0005f",
2488=>x"0005f",
2489=>x"0005f",
2490=>x"0005f",
2491=>x"0005f",
2492=>x"0005f",
2493=>x"0005f",
2494=>x"0005f",
2495=>x"0005f",
2496=>x"0005f",
2497=>x"0005f",
2498=>x"0005f",
2499=>x"0005f",
2500=>x"0005f",
2501=>x"0005f",
2502=>x"0005f",
2503=>x"0005f",
2504=>x"0005f",
2505=>x"0005f",
2506=>x"0005f",
2507=>x"0005f",
2508=>x"0005f",
2509=>x"0005f",
2510=>x"0005f",
2511=>x"0005f",
2512=>x"0005f",
2513=>x"0005f",
2514=>x"0005f",
2515=>x"0005f",
2516=>x"0005f",
2517=>x"0005f",
2518=>x"0005f",
2519=>x"0005f",
2520=>x"0005f",
2521=>x"0005f",
2522=>x"0005f",
2523=>x"0005f",
2524=>x"0005f",
2525=>x"0005f",
2526=>x"0005f",
2527=>x"0005f",
2528=>x"0005f",
2529=>x"0005f",
2530=>x"0005f",
2531=>x"0005f",
2532=>x"0005f",
2533=>x"0005f",
2534=>x"0005f",
2535=>x"0005f",
2536=>x"0005f",
2537=>x"0005f",
2538=>x"0005f",
2539=>x"0005f",
2540=>x"0005f",
2541=>x"0005f",
2542=>x"0005f",
2543=>x"0005f",
2544=>x"0005f",
2545=>x"0005f",
2546=>x"0005f",
2547=>x"0005f",
2548=>x"0005f",
2549=>x"0005f",
2550=>x"0005f",
2551=>x"0005f",
2552=>x"0005f",
2553=>x"0005f",
2554=>x"0005f",
2555=>x"0005f",
2556=>x"0005f",
2557=>x"0005f",
2558=>x"0005f",
2559=>x"0005f",
2560=>x"0005f",
2561=>x"0005f",
2562=>x"0005f",
2563=>x"0005f",
2564=>x"0005f",
2565=>x"0005f",
2566=>x"0005f",
2567=>x"0005f",
2568=>x"0005f",
2569=>x"0005f",
2570=>x"0005f",
2571=>x"0005f",
2572=>x"0005f",
2573=>x"0005f",
2574=>x"0005f",
2575=>x"0005f",
2576=>x"0005f",
2577=>x"0005f",
2578=>x"0005f",
2579=>x"0005f",
2580=>x"0005f",
2581=>x"0005f",
2582=>x"0005f",
2583=>x"0005f",
2584=>x"0005f",
2585=>x"0005f",
2586=>x"0005f",
2587=>x"0005f",
2588=>x"0005f",
2589=>x"0005f",
2590=>x"0005f",
2591=>x"0005f",
2592=>x"0005f",
2593=>x"0005f",
2594=>x"0005f",
2595=>x"0005f",
2596=>x"0005f",
2597=>x"0005f",
2598=>x"0005f",
2599=>x"0005f",
2600=>x"0005f",
2601=>x"0005f",
2602=>x"0005f",
2603=>x"0005f",
2604=>x"0005f",
2605=>x"0005f",
2606=>x"0005f",
2607=>x"0005f",
2608=>x"0005f",
2609=>x"0005f",
2610=>x"0005f",
2611=>x"0005f",
2612=>x"0005f",
2613=>x"0005f",
2614=>x"0005f",
2615=>x"0005f",
2616=>x"0005f",
2617=>x"0005f",
2618=>x"0005f",
2619=>x"0005f",
2620=>x"0005f",
2621=>x"0005f",
2622=>x"0005f",
2623=>x"0005f",
2624=>x"0005f",
2625=>x"0005f",
2626=>x"0005f",
2627=>x"0005f",
2628=>x"0005f",
2629=>x"0005f",
2630=>x"0005f",
2631=>x"0005f",
2632=>x"0005f",
2633=>x"0005f",
2634=>x"0005f",
2635=>x"0005f",
2636=>x"0005f",
2637=>x"0005f",
2638=>x"0005f",
2639=>x"0005f",
2640=>x"0005f",
2641=>x"0005f",
2642=>x"0005f",
2643=>x"0005f",
2644=>x"0005f",
2645=>x"0005f",
2646=>x"0005f",
2647=>x"0005f",
2648=>x"0005f",
2649=>x"0005f",
2650=>x"0005f",
2651=>x"0005f",
2652=>x"0005f",
2653=>x"0005f",
2654=>x"0005f",
2655=>x"0005f",
2656=>x"0005f",
2657=>x"0005f",
2658=>x"0005f",
2659=>x"0005f",
2660=>x"0005f",
2661=>x"0005f",
2662=>x"0005f",
2663=>x"0005f",
2664=>x"0005f",
2665=>x"0005f",
2666=>x"0005f",
2667=>x"0005f",
2668=>x"0005f",
2669=>x"0005f",
2670=>x"0005f",
2671=>x"0005f",
2672=>x"0005f",
2673=>x"0005f",
2674=>x"0005f",
2675=>x"0005f",
2676=>x"0005f",
2677=>x"0005f",
2678=>x"0005f",
2679=>x"0005f",
2680=>x"0005f",
2681=>x"0005f",
2682=>x"0005f",
2683=>x"0005f",
2684=>x"0005f",
2685=>x"0005f",
2686=>x"0005f",
2687=>x"0005f",
2688=>x"0005f",
2689=>x"0005f",
2690=>x"0005f",
2691=>x"0005f",
2692=>x"0005f",
2693=>x"0005f",
2694=>x"0005f",
2695=>x"0005f",
2696=>x"0005f",
2697=>x"0005f",
2698=>x"0005f",
2699=>x"0005f",
2700=>x"0005f",
2701=>x"0005f",
2702=>x"0005f",
2703=>x"0005f",
2704=>x"0005f",
2705=>x"0005f",
2706=>x"0005f",
2707=>x"0005f",
2708=>x"0005f",
2709=>x"0005f",
2710=>x"0005f",
2711=>x"0005f",
2712=>x"0005f",
2713=>x"0005f",
2714=>x"0005f",
2715=>x"0005f",
2716=>x"0005f",
2717=>x"0005f",
2718=>x"0005f",
2719=>x"0005f",
2720=>x"0005f",
2721=>x"0005f",
2722=>x"0005f",
2723=>x"0005f",
2724=>x"0005f",
2725=>x"0005f",
2726=>x"0005f",
2727=>x"0005f",
2728=>x"0005f",
2729=>x"0005f",
2730=>x"0005f",
2731=>x"0005f",
2732=>x"0005f",
2733=>x"0005f",
2734=>x"0005f",
2735=>x"0005f",
2736=>x"0005f",
2737=>x"0005f",
2738=>x"0005f",
2739=>x"0005f",
2740=>x"0005f",
2741=>x"0005f",
2742=>x"0005f",
2743=>x"0005f",
2744=>x"0005f",
2745=>x"0005f",
2746=>x"0005f",
2747=>x"0005f",
2748=>x"0005f",
2749=>x"0005f",
2750=>x"0005f",
2751=>x"0005f",
2752=>x"0005f",
2753=>x"0005f",
2754=>x"0005f",
2755=>x"0005f",
2756=>x"0005f",
2757=>x"0005f",
2758=>x"0005f",
2759=>x"0005f",
2760=>x"0005f",
2761=>x"0005f",
2762=>x"0005f",
2763=>x"0005f",
2764=>x"0005f",
2765=>x"0005f",
2766=>x"0005f",
2767=>x"0005f",
2768=>x"0005f",
2769=>x"0005f",
2770=>x"0005f",
2771=>x"0005f",
2772=>x"0005f",
2773=>x"0005f",
2774=>x"0005f",
2775=>x"0005f",
2776=>x"0005f",
2777=>x"0005f",
2778=>x"0005f",
2779=>x"0005f",
2780=>x"0005f",
2781=>x"0005f",
2782=>x"0005f",
2783=>x"0005f",
2784=>x"0005f",
2785=>x"0005f",
2786=>x"0005f",
2787=>x"0005f",
2788=>x"0005f",
2789=>x"0005f",
2790=>x"0005f",
2791=>x"0005f",
2792=>x"0005f",
2793=>x"0005f",
2794=>x"0005f",
2795=>x"0005f",
2796=>x"0005f",
2797=>x"0005f",
2798=>x"0005f",
2799=>x"0005f",
2800=>x"0005f",
2801=>x"0005f",
2802=>x"0005f",
2803=>x"0005f",
2804=>x"0005f",
2805=>x"0005f",
2806=>x"0005f",
2807=>x"0005f",
2808=>x"0005f",
2809=>x"0005f",
2810=>x"0005f",
2811=>x"0005f",
2812=>x"0005f",
2813=>x"0005f",
2814=>x"0005f",
2815=>x"0005f",
2816=>x"0005f",
2817=>x"0005f",
2818=>x"0005f",
2819=>x"0005f",
2820=>x"0005f",
2821=>x"0005f",
2822=>x"0005f",
2823=>x"0005f",
2824=>x"0005f",
2825=>x"0005f",
2826=>x"0005f",
2827=>x"0005f",
2828=>x"0005f",
2829=>x"0005f",
2830=>x"0005f",
2831=>x"0005f",
2832=>x"0005f",
2833=>x"0005f",
2834=>x"0005f",
2835=>x"0005f",
2836=>x"0005f",
2837=>x"0005f",
2838=>x"0005f",
2839=>x"0005f",
2840=>x"0005f",
2841=>x"0005f",
2842=>x"0005f",
2843=>x"0005f",
2844=>x"0005f",
2845=>x"0005f",
2846=>x"0005f",
2847=>x"0005f",
2848=>x"0005f",
2849=>x"0005f",
2850=>x"0005f",
2851=>x"0005f",
2852=>x"0005f",
2853=>x"0005f",
2854=>x"0005f",
2855=>x"0005f",
2856=>x"0005f",
2857=>x"0005f",
2858=>x"0005f",
2859=>x"0005f",
2860=>x"0005f",
2861=>x"0005f",
2862=>x"0005f",
2863=>x"0005f",
2864=>x"0005f",
2865=>x"0005f",
2866=>x"0005f",
2867=>x"0005f",
2868=>x"0005f",
2869=>x"0005f",
2870=>x"0005f",
2871=>x"0005f",
2872=>x"0005f",
2873=>x"0005f",
2874=>x"0005f",
2875=>x"0005f",
2876=>x"0005f",
2877=>x"0005f",
2878=>x"0005f",
2879=>x"0005f",
2880=>x"0005f",
2881=>x"0005f",
2882=>x"0005f",
2883=>x"0005f",
2884=>x"0005f",
2885=>x"0005f",
2886=>x"0005f",
2887=>x"0005f",
2888=>x"0005f",
2889=>x"0005f",
2890=>x"0005f",
2891=>x"0005f",
2892=>x"0005f",
2893=>x"0005f",
2894=>x"0005f",
2895=>x"0005f",
2896=>x"0005f",
2897=>x"0005f",
2898=>x"0005f",
2899=>x"0005f",
2900=>x"0005f",
2901=>x"0005f",
2902=>x"0005f",
2903=>x"0005f",
2904=>x"0005f",
2905=>x"0005f",
2906=>x"0005f",
2907=>x"0005f",
2908=>x"0005f",
2909=>x"0005f",
2910=>x"0005f",
2911=>x"0005f",
2912=>x"0005f",
2913=>x"0005f",
2914=>x"0005f",
2915=>x"0005f",
2916=>x"0005f",
2917=>x"0005f",
2918=>x"0005f",
2919=>x"0005f",
2920=>x"0005f",
2921=>x"0005f",
2922=>x"0005f",
2923=>x"0005f",
2924=>x"0005f",
2925=>x"0005f",
2926=>x"0005f",
2927=>x"0005f",
2928=>x"0005f",
2929=>x"0005f",
2930=>x"0005f",
2931=>x"0005f",
2932=>x"0005f",
2933=>x"0005f",
2934=>x"0005f",
2935=>x"0005f",
2936=>x"0005f",
2937=>x"0005f",
2938=>x"0005f",
2939=>x"0005f",
2940=>x"0005f",
2941=>x"0005f",
2942=>x"0005f",
2943=>x"0005f",
2944=>x"0005f",
2945=>x"0005f",
2946=>x"0005f",
2947=>x"0005f",
2948=>x"0005f",
2949=>x"0005f",
2950=>x"0005f",
2951=>x"0005f",
2952=>x"0005f",
2953=>x"0005f",
2954=>x"0005f",
2955=>x"0005f",
2956=>x"0005f",
2957=>x"0005f",
2958=>x"0005f",
2959=>x"0005f",
2960=>x"0005f",
2961=>x"0005f",
2962=>x"0005f",
2963=>x"0005f",
2964=>x"0005f",
2965=>x"0005f",
2966=>x"0005f",
2967=>x"0005f",
2968=>x"0005f",
2969=>x"0005f",
2970=>x"0005f",
2971=>x"0005f",
2972=>x"0005f",
2973=>x"0005f",
2974=>x"0005f",
2975=>x"0005f",
2976=>x"0005f",
2977=>x"0005f",
2978=>x"0005f",
2979=>x"0005f",
2980=>x"0005f",
2981=>x"0005f",
2982=>x"0005f",
2983=>x"0005f",
2984=>x"0005f",
2985=>x"0005f",
2986=>x"0005f",
2987=>x"0005f",
2988=>x"0005f",
2989=>x"0005f",
2990=>x"0005f",
2991=>x"0005f",
2992=>x"0005f",
2993=>x"0005f",
2994=>x"0005f",
2995=>x"0005f",
2996=>x"0005f",
2997=>x"0005f",
2998=>x"0005f",
2999=>x"0005f",
3000=>x"0005f",
3001=>x"0005f",
3002=>x"0005f",
3003=>x"0005f",
3004=>x"0005f",
3005=>x"0005f",
3006=>x"0005f",
3007=>x"0005f",
3008=>x"0005f",
3009=>x"0005f",
3010=>x"0005f",
3011=>x"0005f",
3012=>x"0005f",
3013=>x"0005f",
3014=>x"0005f",
3015=>x"0005f",
3016=>x"0005f",
3017=>x"0005f",
3018=>x"0005f",
3019=>x"0005f",
3020=>x"0005f",
3021=>x"0005f",
3022=>x"0005f",
3023=>x"0005f",
3024=>x"0005f",
3025=>x"0005f",
3026=>x"0005f",
3027=>x"0005f",
3028=>x"0005f",
3029=>x"0005f",
3030=>x"0005f",
3031=>x"0005f",
3032=>x"0005f",
3033=>x"0005f",
3034=>x"0005f",
3035=>x"0005f",
3036=>x"0005f",
3037=>x"0005f",
3038=>x"0005f",
3039=>x"0005f",
3040=>x"0005f",
3041=>x"0005f",
3042=>x"0005f",
3043=>x"0005f",
3044=>x"0005f",
3045=>x"0005f",
3046=>x"0005f",
3047=>x"0005f",
3048=>x"0005f",
3049=>x"0005f",
3050=>x"0005f",
3051=>x"0005f",
3052=>x"0005f",
3053=>x"0005f",
3054=>x"0005f",
3055=>x"0005f",
3056=>x"0005f",
3057=>x"0005f",
3058=>x"0005f",
3059=>x"0005f",
3060=>x"0005f",
3061=>x"0005f",
3062=>x"0005f",
3063=>x"0005f",
3064=>x"0005f",
3065=>x"0005f",
3066=>x"0005f",
3067=>x"0005f",
3068=>x"0005f",
3069=>x"0005f",
3070=>x"0005f",
3071=>x"0005f",
3072=>x"00060",
3073=>x"00060",
3074=>x"00060",
3075=>x"00060",
3076=>x"00060",
3077=>x"00060",
3078=>x"00060",
3079=>x"00060",
3080=>x"00060",
3081=>x"00060",
3082=>x"00060",
3083=>x"00060",
3084=>x"00060",
3085=>x"00060",
3086=>x"00060",
3087=>x"00060",
3088=>x"00060",
3089=>x"00060",
3090=>x"00060",
3091=>x"00060",
3092=>x"00060",
3093=>x"00060",
3094=>x"00060",
3095=>x"00060",
3096=>x"00060",
3097=>x"00060",
3098=>x"00060",
3099=>x"00060",
3100=>x"00060",
3101=>x"00060",
3102=>x"00060",
3103=>x"00060",
3104=>x"00060",
3105=>x"00060",
3106=>x"00060",
3107=>x"00060",
3108=>x"00060",
3109=>x"00060",
3110=>x"00060",
3111=>x"00060",
3112=>x"00060",
3113=>x"00060",
3114=>x"00060",
3115=>x"00060",
3116=>x"00060",
3117=>x"00060",
3118=>x"00060",
3119=>x"00060",
3120=>x"00060",
3121=>x"00060",
3122=>x"00060",
3123=>x"00060",
3124=>x"00060",
3125=>x"00060",
3126=>x"00060",
3127=>x"00060",
3128=>x"00060",
3129=>x"00060",
3130=>x"00060",
3131=>x"00060",
3132=>x"00060",
3133=>x"00060",
3134=>x"00060",
3135=>x"00060",
3136=>x"00060",
3137=>x"00060",
3138=>x"00060",
3139=>x"00060",
3140=>x"00060",
3141=>x"00060",
3142=>x"00060",
3143=>x"00060",
3144=>x"00060",
3145=>x"00060",
3146=>x"00060",
3147=>x"00060",
3148=>x"00060",
3149=>x"00060",
3150=>x"00060",
3151=>x"00060",
3152=>x"00060",
3153=>x"00060",
3154=>x"00060",
3155=>x"00060",
3156=>x"00060",
3157=>x"00060",
3158=>x"00060",
3159=>x"00060",
3160=>x"00060",
3161=>x"00060",
3162=>x"00060",
3163=>x"00060",
3164=>x"00060",
3165=>x"00060",
3166=>x"00060",
3167=>x"00060",
3168=>x"00060",
3169=>x"00060",
3170=>x"00060",
3171=>x"00060",
3172=>x"00060",
3173=>x"00060",
3174=>x"00060",
3175=>x"00060",
3176=>x"00060",
3177=>x"00060",
3178=>x"00060",
3179=>x"00060",
3180=>x"00060",
3181=>x"00060",
3182=>x"00060",
3183=>x"00060",
3184=>x"00060",
3185=>x"00060",
3186=>x"00060",
3187=>x"00060",
3188=>x"00060",
3189=>x"00060",
3190=>x"00060",
3191=>x"00060",
3192=>x"00060",
3193=>x"00060",
3194=>x"00060",
3195=>x"00060",
3196=>x"00060",
3197=>x"00060",
3198=>x"00060",
3199=>x"00060",
3200=>x"00060",
3201=>x"00060",
3202=>x"00060",
3203=>x"00060",
3204=>x"00060",
3205=>x"00060",
3206=>x"00060",
3207=>x"00060",
3208=>x"00060",
3209=>x"00060",
3210=>x"00060",
3211=>x"00060",
3212=>x"00060",
3213=>x"00060",
3214=>x"00060",
3215=>x"00060",
3216=>x"00060",
3217=>x"00060",
3218=>x"00060",
3219=>x"00060",
3220=>x"00060",
3221=>x"00060",
3222=>x"00060",
3223=>x"00060",
3224=>x"00060",
3225=>x"00060",
3226=>x"00060",
3227=>x"00060",
3228=>x"00060",
3229=>x"00060",
3230=>x"00060",
3231=>x"00060",
3232=>x"00060",
3233=>x"00060",
3234=>x"00060",
3235=>x"00060",
3236=>x"00060",
3237=>x"00060",
3238=>x"00060",
3239=>x"00060",
3240=>x"00060",
3241=>x"00060",
3242=>x"00060",
3243=>x"00060",
3244=>x"00060",
3245=>x"00060",
3246=>x"00060",
3247=>x"00060",
3248=>x"00060",
3249=>x"00060",
3250=>x"00060",
3251=>x"00060",
3252=>x"00060",
3253=>x"00060",
3254=>x"00060",
3255=>x"00060",
3256=>x"00060",
3257=>x"00060",
3258=>x"00060",
3259=>x"00060",
3260=>x"00060",
3261=>x"00060",
3262=>x"00060",
3263=>x"00060",
3264=>x"00060",
3265=>x"00060",
3266=>x"00060",
3267=>x"00060",
3268=>x"00060",
3269=>x"00060",
3270=>x"00060",
3271=>x"00060",
3272=>x"00060",
3273=>x"00060",
3274=>x"00060",
3275=>x"00060",
3276=>x"00060",
3277=>x"00060",
3278=>x"00060",
3279=>x"00060",
3280=>x"00060",
3281=>x"00060",
3282=>x"00060",
3283=>x"00060",
3284=>x"00060",
3285=>x"00060",
3286=>x"00060",
3287=>x"00060",
3288=>x"00060",
3289=>x"00060",
3290=>x"00060",
3291=>x"00060",
3292=>x"00060",
3293=>x"00060",
3294=>x"00060",
3295=>x"00060",
3296=>x"00060",
3297=>x"00060",
3298=>x"00060",
3299=>x"00060",
3300=>x"00060",
3301=>x"00060",
3302=>x"00060",
3303=>x"00060",
3304=>x"00060",
3305=>x"00060",
3306=>x"00060",
3307=>x"00060",
3308=>x"00060",
3309=>x"00060",
3310=>x"00060",
3311=>x"00060",
3312=>x"00060",
3313=>x"00060",
3314=>x"00060",
3315=>x"00060",
3316=>x"00060",
3317=>x"00060",
3318=>x"00060",
3319=>x"00060",
3320=>x"00060",
3321=>x"00060",
3322=>x"00060",
3323=>x"00060",
3324=>x"00060",
3325=>x"00060",
3326=>x"00060",
3327=>x"00060",
3328=>x"00060",
3329=>x"00060",
3330=>x"00060",
3331=>x"00060",
3332=>x"00060",
3333=>x"00060",
3334=>x"00060",
3335=>x"00060",
3336=>x"00060",
3337=>x"00060",
3338=>x"00060",
3339=>x"00060",
3340=>x"00060",
3341=>x"00060",
3342=>x"00060",
3343=>x"00060",
3344=>x"00060",
3345=>x"00060",
3346=>x"00060",
3347=>x"00060",
3348=>x"00060",
3349=>x"00060",
3350=>x"00060",
3351=>x"00060",
3352=>x"00060",
3353=>x"00060",
3354=>x"00060",
3355=>x"00060",
3356=>x"00060",
3357=>x"00060",
3358=>x"00060",
3359=>x"00060",
3360=>x"00060",
3361=>x"00060",
3362=>x"00060",
3363=>x"00060",
3364=>x"00060",
3365=>x"00060",
3366=>x"00060",
3367=>x"00060",
3368=>x"00060",
3369=>x"00060",
3370=>x"00060",
3371=>x"00060",
3372=>x"00060",
3373=>x"00060",
3374=>x"00060",
3375=>x"00060",
3376=>x"00060",
3377=>x"00060",
3378=>x"00060",
3379=>x"00060",
3380=>x"00060",
3381=>x"00060",
3382=>x"00060",
3383=>x"00060",
3384=>x"00060",
3385=>x"00060",
3386=>x"00060",
3387=>x"00060",
3388=>x"00060",
3389=>x"00060",
3390=>x"00060",
3391=>x"00060",
3392=>x"00060",
3393=>x"00060",
3394=>x"00060",
3395=>x"00060",
3396=>x"00060",
3397=>x"00060",
3398=>x"00060",
3399=>x"00060",
3400=>x"00060",
3401=>x"00060",
3402=>x"00060",
3403=>x"00060",
3404=>x"00060",
3405=>x"00060",
3406=>x"00060",
3407=>x"00060",
3408=>x"00060",
3409=>x"00060",
3410=>x"00060",
3411=>x"00060",
3412=>x"00060",
3413=>x"00060",
3414=>x"00060",
3415=>x"00060",
3416=>x"00060",
3417=>x"00060",
3418=>x"00060",
3419=>x"00060",
3420=>x"00060",
3421=>x"00060",
3422=>x"00060",
3423=>x"00060",
3424=>x"00060",
3425=>x"00060",
3426=>x"00060",
3427=>x"00060",
3428=>x"00060",
3429=>x"00060",
3430=>x"00060",
3431=>x"00060",
3432=>x"00060",
3433=>x"00060",
3434=>x"00060",
3435=>x"00060",
3436=>x"00060",
3437=>x"00060",
3438=>x"00060",
3439=>x"00060",
3440=>x"00060",
3441=>x"00060",
3442=>x"00060",
3443=>x"00060",
3444=>x"00060",
3445=>x"00060",
3446=>x"00060",
3447=>x"00060",
3448=>x"00060",
3449=>x"00060",
3450=>x"00060",
3451=>x"00060",
3452=>x"00060",
3453=>x"00060",
3454=>x"00060",
3455=>x"00060",
3456=>x"00060",
3457=>x"00060",
3458=>x"00060",
3459=>x"00060",
3460=>x"00060",
3461=>x"00060",
3462=>x"00060",
3463=>x"00060",
3464=>x"00060",
3465=>x"00060",
3466=>x"00060",
3467=>x"00060",
3468=>x"00060",
3469=>x"00060",
3470=>x"00060",
3471=>x"00060",
3472=>x"00060",
3473=>x"00060",
3474=>x"00060",
3475=>x"00060",
3476=>x"00060",
3477=>x"00060",
3478=>x"00060",
3479=>x"00060",
3480=>x"00060",
3481=>x"00060",
3482=>x"00060",
3483=>x"00060",
3484=>x"00060",
3485=>x"00060",
3486=>x"00060",
3487=>x"00060",
3488=>x"00060",
3489=>x"00060",
3490=>x"00060",
3491=>x"00060",
3492=>x"00060",
3493=>x"00060",
3494=>x"00060",
3495=>x"00060",
3496=>x"00060",
3497=>x"00060",
3498=>x"00060",
3499=>x"00060",
3500=>x"00060",
3501=>x"00060",
3502=>x"00060",
3503=>x"00060",
3504=>x"00060",
3505=>x"00060",
3506=>x"00060",
3507=>x"00060",
3508=>x"00060",
3509=>x"00060",
3510=>x"00060",
3511=>x"00060",
3512=>x"00060",
3513=>x"00060",
3514=>x"00060",
3515=>x"00060",
3516=>x"00060",
3517=>x"00060",
3518=>x"00060",
3519=>x"00060",
3520=>x"00060",
3521=>x"00060",
3522=>x"00060",
3523=>x"00060",
3524=>x"00060",
3525=>x"00060",
3526=>x"00060",
3527=>x"00060",
3528=>x"00060",
3529=>x"00060",
3530=>x"00060",
3531=>x"00060",
3532=>x"00060",
3533=>x"00060",
3534=>x"00060",
3535=>x"00060",
3536=>x"00060",
3537=>x"00060",
3538=>x"00060",
3539=>x"00060",
3540=>x"00060",
3541=>x"00060",
3542=>x"00060",
3543=>x"00060",
3544=>x"00060",
3545=>x"00060",
3546=>x"00060",
3547=>x"00060",
3548=>x"00060",
3549=>x"00060",
3550=>x"00060",
3551=>x"00060",
3552=>x"00060",
3553=>x"00060",
3554=>x"00060",
3555=>x"00060",
3556=>x"00060",
3557=>x"00060",
3558=>x"00060",
3559=>x"00060",
3560=>x"00060",
3561=>x"00060",
3562=>x"00060",
3563=>x"00060",
3564=>x"00060",
3565=>x"00060",
3566=>x"00060",
3567=>x"00060",
3568=>x"00060",
3569=>x"00060",
3570=>x"00060",
3571=>x"00060",
3572=>x"00060",
3573=>x"00060",
3574=>x"00060",
3575=>x"00060",
3576=>x"00060",
3577=>x"00060",
3578=>x"00060",
3579=>x"00060",
3580=>x"00060",
3581=>x"00060",
3582=>x"00060",
3583=>x"00060",
3584=>x"00060",
3585=>x"00060",
3586=>x"00060",
3587=>x"00060",
3588=>x"00060",
3589=>x"00060",
3590=>x"00060",
3591=>x"00060",
3592=>x"00060",
3593=>x"00060",
3594=>x"00060",
3595=>x"00060",
3596=>x"00060",
3597=>x"00060",
3598=>x"00060",
3599=>x"00060",
3600=>x"00060",
3601=>x"00060",
3602=>x"00060",
3603=>x"00060",
3604=>x"00060",
3605=>x"00060",
3606=>x"00060",
3607=>x"00060",
3608=>x"00060",
3609=>x"00060",
3610=>x"00060",
3611=>x"00060",
3612=>x"00060",
3613=>x"00060",
3614=>x"00060",
3615=>x"00060",
3616=>x"00060",
3617=>x"00060",
3618=>x"00060",
3619=>x"00060",
3620=>x"00060",
3621=>x"00060",
3622=>x"00060",
3623=>x"00060",
3624=>x"00060",
3625=>x"00060",
3626=>x"00060",
3627=>x"00060",
3628=>x"00060",
3629=>x"00060",
3630=>x"00060",
3631=>x"00060",
3632=>x"00060",
3633=>x"00060",
3634=>x"00060",
3635=>x"00060",
3636=>x"00060",
3637=>x"00060",
3638=>x"00060",
3639=>x"00060",
3640=>x"00060",
3641=>x"00060",
3642=>x"00060",
3643=>x"00060",
3644=>x"00060",
3645=>x"00060",
3646=>x"00060",
3647=>x"00060",
3648=>x"00060",
3649=>x"00060",
3650=>x"00060",
3651=>x"00060",
3652=>x"00060",
3653=>x"00060",
3654=>x"00060",
3655=>x"00060",
3656=>x"00060",
3657=>x"00060",
3658=>x"00060",
3659=>x"00060",
3660=>x"00060",
3661=>x"00060",
3662=>x"00060",
3663=>x"00060",
3664=>x"00060",
3665=>x"00060",
3666=>x"00060",
3667=>x"00060",
3668=>x"00060",
3669=>x"00060",
3670=>x"00060",
3671=>x"00060",
3672=>x"00060",
3673=>x"00060",
3674=>x"00060",
3675=>x"00060",
3676=>x"00060",
3677=>x"00060",
3678=>x"00060",
3679=>x"00060",
3680=>x"00060",
3681=>x"00060",
3682=>x"00060",
3683=>x"00060",
3684=>x"00060",
3685=>x"00060",
3686=>x"00060",
3687=>x"00060",
3688=>x"00060",
3689=>x"00060",
3690=>x"00060",
3691=>x"00060",
3692=>x"00060",
3693=>x"00060",
3694=>x"00060",
3695=>x"00060",
3696=>x"00060",
3697=>x"00060",
3698=>x"00060",
3699=>x"00060",
3700=>x"00060",
3701=>x"00060",
3702=>x"00060",
3703=>x"00060",
3704=>x"00060",
3705=>x"00060",
3706=>x"00060",
3707=>x"00060",
3708=>x"00060",
3709=>x"00060",
3710=>x"00060",
3711=>x"00060",
3712=>x"00060",
3713=>x"00060",
3714=>x"00060",
3715=>x"00060",
3716=>x"00060",
3717=>x"00060",
3718=>x"00060",
3719=>x"00060",
3720=>x"00060",
3721=>x"00060",
3722=>x"00060",
3723=>x"00060",
3724=>x"00060",
3725=>x"00060",
3726=>x"00060",
3727=>x"00060",
3728=>x"00060",
3729=>x"00060",
3730=>x"00060",
3731=>x"00060",
3732=>x"00060",
3733=>x"00060",
3734=>x"00060",
3735=>x"00060",
3736=>x"00060",
3737=>x"00060",
3738=>x"00060",
3739=>x"00060",
3740=>x"00060",
3741=>x"00060",
3742=>x"00060",
3743=>x"00060",
3744=>x"00060",
3745=>x"00060",
3746=>x"00060",
3747=>x"00060",
3748=>x"00060",
3749=>x"00060",
3750=>x"00060",
3751=>x"00060",
3752=>x"00060",
3753=>x"00060",
3754=>x"00060",
3755=>x"00060",
3756=>x"00060",
3757=>x"00060",
3758=>x"00060",
3759=>x"00060",
3760=>x"00060",
3761=>x"00060",
3762=>x"00060",
3763=>x"00060",
3764=>x"00060",
3765=>x"00060",
3766=>x"00060",
3767=>x"00060",
3768=>x"00060",
3769=>x"00060",
3770=>x"00060",
3771=>x"00060",
3772=>x"00060",
3773=>x"00060",
3774=>x"00060",
3775=>x"00060",
3776=>x"00060",
3777=>x"00060",
3778=>x"00060",
3779=>x"00060",
3780=>x"00060",
3781=>x"00060",
3782=>x"00060",
3783=>x"00060",
3784=>x"00060",
3785=>x"00060",
3786=>x"00060",
3787=>x"00060",
3788=>x"00060",
3789=>x"00060",
3790=>x"00060",
3791=>x"00060",
3792=>x"00060",
3793=>x"00060",
3794=>x"00060",
3795=>x"00060",
3796=>x"00060",
3797=>x"00060",
3798=>x"00060",
3799=>x"00060",
3800=>x"00060",
3801=>x"00060",
3802=>x"00060",
3803=>x"00060",
3804=>x"00060",
3805=>x"00060",
3806=>x"00060",
3807=>x"00060",
3808=>x"00060",
3809=>x"00060",
3810=>x"00060",
3811=>x"00060",
3812=>x"00060",
3813=>x"00060",
3814=>x"00060",
3815=>x"00060",
3816=>x"00060",
3817=>x"00060",
3818=>x"00060",
3819=>x"00060",
3820=>x"00060",
3821=>x"00060",
3822=>x"00060",
3823=>x"00060",
3824=>x"00060",
3825=>x"00060",
3826=>x"00060",
3827=>x"00060",
3828=>x"00060",
3829=>x"00060",
3830=>x"00060",
3831=>x"00060",
3832=>x"00060",
3833=>x"00060",
3834=>x"00060",
3835=>x"00060",
3836=>x"00060",
3837=>x"00060",
3838=>x"00060",
3839=>x"00060",
3840=>x"00060",
3841=>x"00060",
3842=>x"00060",
3843=>x"00060",
3844=>x"00060",
3845=>x"00060",
3846=>x"00060",
3847=>x"00060",
3848=>x"00060",
3849=>x"00060",
3850=>x"00060",
3851=>x"00060",
3852=>x"00060",
3853=>x"00060",
3854=>x"00060",
3855=>x"00060",
3856=>x"00060",
3857=>x"00060",
3858=>x"00060",
3859=>x"00060",
3860=>x"00060",
3861=>x"00060",
3862=>x"00060",
3863=>x"00060",
3864=>x"00060",
3865=>x"00060",
3866=>x"00060",
3867=>x"00060",
3868=>x"00060",
3869=>x"00060",
3870=>x"00060",
3871=>x"00060",
3872=>x"00060",
3873=>x"00060",
3874=>x"00060",
3875=>x"00060",
3876=>x"00060",
3877=>x"00060",
3878=>x"00060",
3879=>x"00060",
3880=>x"00060",
3881=>x"00060",
3882=>x"00060",
3883=>x"00060",
3884=>x"00060",
3885=>x"00060",
3886=>x"00060",
3887=>x"00060",
3888=>x"00060",
3889=>x"00060",
3890=>x"00060",
3891=>x"00060",
3892=>x"00060",
3893=>x"00060",
3894=>x"00060",
3895=>x"00060",
3896=>x"00060",
3897=>x"00060",
3898=>x"00060",
3899=>x"00060",
3900=>x"00060",
3901=>x"00060",
3902=>x"00060",
3903=>x"00060",
3904=>x"00060",
3905=>x"00060",
3906=>x"00060",
3907=>x"00060",
3908=>x"00060",
3909=>x"00060",
3910=>x"00060",
3911=>x"00060",
3912=>x"00060",
3913=>x"00060",
3914=>x"00060",
3915=>x"00060",
3916=>x"00060",
3917=>x"00060",
3918=>x"00060",
3919=>x"00060",
3920=>x"00060",
3921=>x"00060",
3922=>x"00060",
3923=>x"00060",
3924=>x"00060",
3925=>x"00060",
3926=>x"00060",
3927=>x"00060",
3928=>x"00060",
3929=>x"00060",
3930=>x"00060",
3931=>x"00060",
3932=>x"00060",
3933=>x"00060",
3934=>x"00060",
3935=>x"00060",
3936=>x"00060",
3937=>x"00060",
3938=>x"00060",
3939=>x"00060",
3940=>x"00060",
3941=>x"00060",
3942=>x"00060",
3943=>x"00060",
3944=>x"00060",
3945=>x"00060",
3946=>x"00060",
3947=>x"00060",
3948=>x"00060",
3949=>x"00060",
3950=>x"00060",
3951=>x"00060",
3952=>x"00060",
3953=>x"00060",
3954=>x"00060",
3955=>x"00060",
3956=>x"00060",
3957=>x"00060",
3958=>x"00060",
3959=>x"00060",
3960=>x"00060",
3961=>x"00060",
3962=>x"00060",
3963=>x"00060",
3964=>x"00060",
3965=>x"00060",
3966=>x"00060",
3967=>x"00060",
3968=>x"00060",
3969=>x"00060",
3970=>x"00060",
3971=>x"00060",
3972=>x"00060",
3973=>x"00060",
3974=>x"00060",
3975=>x"00060",
3976=>x"00060",
3977=>x"00060",
3978=>x"00060",
3979=>x"00060",
3980=>x"00060",
3981=>x"00060",
3982=>x"00060",
3983=>x"00060",
3984=>x"00060",
3985=>x"00060",
3986=>x"00060",
3987=>x"00060",
3988=>x"00060",
3989=>x"00060",
3990=>x"00060",
3991=>x"00060",
3992=>x"00060",
3993=>x"00060",
3994=>x"00060",
3995=>x"00060",
3996=>x"00060",
3997=>x"00060",
3998=>x"00060",
3999=>x"00060",
4000=>x"00060",
4001=>x"00060",
4002=>x"00060",
4003=>x"00060",
4004=>x"00060",
4005=>x"00060",
4006=>x"00060",
4007=>x"00060",
4008=>x"00060",
4009=>x"00060",
4010=>x"00060",
4011=>x"00060",
4012=>x"00060",
4013=>x"00060",
4014=>x"00060",
4015=>x"00060",
4016=>x"00060",
4017=>x"00060",
4018=>x"00060",
4019=>x"00060",
4020=>x"00060",
4021=>x"00060",
4022=>x"00060",
4023=>x"00060",
4024=>x"00060",
4025=>x"00060",
4026=>x"00060",
4027=>x"00060",
4028=>x"00060",
4029=>x"00060",
4030=>x"00060",
4031=>x"00060",
4032=>x"00060",
4033=>x"00060",
4034=>x"00060",
4035=>x"00060",
4036=>x"00060",
4037=>x"00060",
4038=>x"00060",
4039=>x"00060",
4040=>x"00060",
4041=>x"00060",
4042=>x"00060",
4043=>x"00060",
4044=>x"00060",
4045=>x"00060",
4046=>x"00060",
4047=>x"00060",
4048=>x"00060",
4049=>x"00060",
4050=>x"00060",
4051=>x"00060",
4052=>x"00060",
4053=>x"00060",
4054=>x"00060",
4055=>x"00060",
4056=>x"00060",
4057=>x"00060",
4058=>x"00060",
4059=>x"00060",
4060=>x"00060",
4061=>x"00060",
4062=>x"00060",
4063=>x"00060",
4064=>x"00060",
4065=>x"00060",
4066=>x"00060",
4067=>x"00060",
4068=>x"00060",
4069=>x"00060",
4070=>x"00060",
4071=>x"00060",
4072=>x"00060",
4073=>x"00060",
4074=>x"00060",
4075=>x"00060",
4076=>x"00060",
4077=>x"00060",
4078=>x"00060",
4079=>x"00060",
4080=>x"00060",
4081=>x"00060",
4082=>x"00060",
4083=>x"00060",
4084=>x"00060",
4085=>x"00060",
4086=>x"00060",
4087=>x"00060",
4088=>x"00060",
4089=>x"00060",
4090=>x"00060",
4091=>x"00060",
4092=>x"00060",
4093=>x"00060",
4094=>x"00060",

others=>x"00000"
);
begin
Cout<=memory(to_integer(unsigned(addr)));

end Behavioral;
