library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.ALL;

entity RSI_ROM2 is
    Port ( addr : in STD_LOGIC_VECTOR (11 downto 0);
           Cout : out STD_LOGIC_VECTOR (19 downto 0));
end RSI_ROM2;

architecture Behavioral of RSI_ROM2 is
type vector is Array(0 to 4095) of Std_logic_vector(19 downto 0);
Constant memory: vector:=
(
0=>x"00001",
1=>x"00001",
2=>x"00002",
3=>x"00003",
4=>x"00004",
5=>x"00004",
6=>x"00005",
7=>x"00006",
8=>x"00006",
9=>x"00007",
10=>x"00008",
11=>x"00008",
12=>x"00009",
13=>x"0000a",
14=>x"0000a",
15=>x"0000b",
16=>x"0000c",
17=>x"0000c",
18=>x"0000d",
19=>x"0000d",
20=>x"0000e",
21=>x"0000f",
22=>x"0000f",
23=>x"00010",
24=>x"00010",
25=>x"00011",
26=>x"00011",
27=>x"00012",
28=>x"00012",
29=>x"00013",
30=>x"00013",
31=>x"00014",
32=>x"00015",
33=>x"00015",
34=>x"00015",
35=>x"00016",
36=>x"00016",
37=>x"00017",
38=>x"00017",
39=>x"00018",
40=>x"00018",
41=>x"00019",
42=>x"00019",
43=>x"0001a",
44=>x"0001a",
45=>x"0001b",
46=>x"0001b",
47=>x"0001b",
48=>x"0001c",
49=>x"0001c",
50=>x"0001d",
51=>x"0001d",
52=>x"0001d",
53=>x"0001e",
54=>x"0001e",
55=>x"0001f",
56=>x"0001f",
57=>x"0001f",
58=>x"00020",
59=>x"00020",
60=>x"00020",
61=>x"00021",
62=>x"00021",
63=>x"00021",
64=>x"00022",
65=>x"00022",
66=>x"00023",
67=>x"00023",
68=>x"00023",
69=>x"00024",
70=>x"00024",
71=>x"00024",
72=>x"00025",
73=>x"00025",
74=>x"00025",
75=>x"00025",
76=>x"00026",
77=>x"00026",
78=>x"00026",
79=>x"00027",
80=>x"00027",
81=>x"00027",
82=>x"00028",
83=>x"00028",
84=>x"00028",
85=>x"00028",
86=>x"00029",
87=>x"00029",
88=>x"00029",
89=>x"0002a",
90=>x"0002a",
91=>x"0002a",
92=>x"0002a",
93=>x"0002b",
94=>x"0002b",
95=>x"0002b",
96=>x"0002b",
97=>x"0002c",
98=>x"0002c",
99=>x"0002c",
100=>x"0002c",
101=>x"0002d",
102=>x"0002d",
103=>x"0002d",
104=>x"0002d",
105=>x"0002e",
106=>x"0002e",
107=>x"0002e",
108=>x"0002e",
109=>x"0002e",
110=>x"0002f",
111=>x"0002f",
112=>x"0002f",
113=>x"0002f",
114=>x"00030",
115=>x"00030",
116=>x"00030",
117=>x"00030",
118=>x"00030",
119=>x"00031",
120=>x"00031",
121=>x"00031",
122=>x"00031",
123=>x"00032",
124=>x"00032",
125=>x"00032",
126=>x"00032",
127=>x"00032",
128=>x"00033",
129=>x"00033",
130=>x"00033",
131=>x"00033",
132=>x"00033",
133=>x"00033",
134=>x"00034",
135=>x"00034",
136=>x"00034",
137=>x"00034",
138=>x"00034",
139=>x"00035",
140=>x"00035",
141=>x"00035",
142=>x"00035",
143=>x"00035",
144=>x"00035",
145=>x"00036",
146=>x"00036",
147=>x"00036",
148=>x"00036",
149=>x"00036",
150=>x"00036",
151=>x"00037",
152=>x"00037",
153=>x"00037",
154=>x"00037",
155=>x"00037",
156=>x"00037",
157=>x"00038",
158=>x"00038",
159=>x"00038",
160=>x"00038",
161=>x"00038",
162=>x"00038",
163=>x"00039",
164=>x"00039",
165=>x"00039",
166=>x"00039",
167=>x"00039",
168=>x"00039",
169=>x"00039",
170=>x"0003a",
171=>x"0003a",
172=>x"0003a",
173=>x"0003a",
174=>x"0003a",
175=>x"0003a",
176=>x"0003a",
177=>x"0003b",
178=>x"0003b",
179=>x"0003b",
180=>x"0003b",
181=>x"0003b",
182=>x"0003b",
183=>x"0003b",
184=>x"0003b",
185=>x"0003c",
186=>x"0003c",
187=>x"0003c",
188=>x"0003c",
189=>x"0003c",
190=>x"0003c",
191=>x"0003c",
192=>x"0003d",
193=>x"0003d",
194=>x"0003d",
195=>x"0003d",
196=>x"0003d",
197=>x"0003d",
198=>x"0003d",
199=>x"0003d",
200=>x"0003d",
201=>x"0003e",
202=>x"0003e",
203=>x"0003e",
204=>x"0003e",
205=>x"0003e",
206=>x"0003e",
207=>x"0003e",
208=>x"0003e",
209=>x"0003f",
210=>x"0003f",
211=>x"0003f",
212=>x"0003f",
213=>x"0003f",
214=>x"0003f",
215=>x"0003f",
216=>x"0003f",
217=>x"0003f",
218=>x"00040",
219=>x"00040",
220=>x"00040",
221=>x"00040",
222=>x"00040",
223=>x"00040",
224=>x"00040",
225=>x"00040",
226=>x"00040",
227=>x"00040",
228=>x"00041",
229=>x"00041",
230=>x"00041",
231=>x"00041",
232=>x"00041",
233=>x"00041",
234=>x"00041",
235=>x"00041",
236=>x"00041",
237=>x"00041",
238=>x"00042",
239=>x"00042",
240=>x"00042",
241=>x"00042",
242=>x"00042",
243=>x"00042",
244=>x"00042",
245=>x"00042",
246=>x"00042",
247=>x"00042",
248=>x"00042",
249=>x"00043",
250=>x"00043",
251=>x"00043",
252=>x"00043",
253=>x"00043",
254=>x"00043",
255=>x"00043",
256=>x"00043",
257=>x"00043",
258=>x"00043",
259=>x"00043",
260=>x"00044",
261=>x"00044",
262=>x"00044",
263=>x"00044",
264=>x"00044",
265=>x"00044",
266=>x"00044",
267=>x"00044",
268=>x"00044",
269=>x"00044",
270=>x"00044",
271=>x"00044",
272=>x"00045",
273=>x"00045",
274=>x"00045",
275=>x"00045",
276=>x"00045",
277=>x"00045",
278=>x"00045",
279=>x"00045",
280=>x"00045",
281=>x"00045",
282=>x"00045",
283=>x"00045",
284=>x"00045",
285=>x"00046",
286=>x"00046",
287=>x"00046",
288=>x"00046",
289=>x"00046",
290=>x"00046",
291=>x"00046",
292=>x"00046",
293=>x"00046",
294=>x"00046",
295=>x"00046",
296=>x"00046",
297=>x"00046",
298=>x"00046",
299=>x"00047",
300=>x"00047",
301=>x"00047",
302=>x"00047",
303=>x"00047",
304=>x"00047",
305=>x"00047",
306=>x"00047",
307=>x"00047",
308=>x"00047",
309=>x"00047",
310=>x"00047",
311=>x"00047",
312=>x"00047",
313=>x"00047",
314=>x"00048",
315=>x"00048",
316=>x"00048",
317=>x"00048",
318=>x"00048",
319=>x"00048",
320=>x"00048",
321=>x"00048",
322=>x"00048",
323=>x"00048",
324=>x"00048",
325=>x"00048",
326=>x"00048",
327=>x"00048",
328=>x"00048",
329=>x"00048",
330=>x"00049",
331=>x"00049",
332=>x"00049",
333=>x"00049",
334=>x"00049",
335=>x"00049",
336=>x"00049",
337=>x"00049",
338=>x"00049",
339=>x"00049",
340=>x"00049",
341=>x"00049",
342=>x"00049",
343=>x"00049",
344=>x"00049",
345=>x"00049",
346=>x"00049",
347=>x"0004a",
348=>x"0004a",
349=>x"0004a",
350=>x"0004a",
351=>x"0004a",
352=>x"0004a",
353=>x"0004a",
354=>x"0004a",
355=>x"0004a",
356=>x"0004a",
357=>x"0004a",
358=>x"0004a",
359=>x"0004a",
360=>x"0004a",
361=>x"0004a",
362=>x"0004a",
363=>x"0004a",
364=>x"0004a",
365=>x"0004b",
366=>x"0004b",
367=>x"0004b",
368=>x"0004b",
369=>x"0004b",
370=>x"0004b",
371=>x"0004b",
372=>x"0004b",
373=>x"0004b",
374=>x"0004b",
375=>x"0004b",
376=>x"0004b",
377=>x"0004b",
378=>x"0004b",
379=>x"0004b",
380=>x"0004b",
381=>x"0004b",
382=>x"0004b",
383=>x"0004b",
384=>x"0004c",
385=>x"0004c",
386=>x"0004c",
387=>x"0004c",
388=>x"0004c",
389=>x"0004c",
390=>x"0004c",
391=>x"0004c",
392=>x"0004c",
393=>x"0004c",
394=>x"0004c",
395=>x"0004c",
396=>x"0004c",
397=>x"0004c",
398=>x"0004c",
399=>x"0004c",
400=>x"0004c",
401=>x"0004c",
402=>x"0004c",
403=>x"0004c",
404=>x"0004c",
405=>x"0004c",
406=>x"0004d",
407=>x"0004d",
408=>x"0004d",
409=>x"0004d",
410=>x"0004d",
411=>x"0004d",
412=>x"0004d",
413=>x"0004d",
414=>x"0004d",
415=>x"0004d",
416=>x"0004d",
417=>x"0004d",
418=>x"0004d",
419=>x"0004d",
420=>x"0004d",
421=>x"0004d",
422=>x"0004d",
423=>x"0004d",
424=>x"0004d",
425=>x"0004d",
426=>x"0004d",
427=>x"0004d",
428=>x"0004d",
429=>x"0004e",
430=>x"0004e",
431=>x"0004e",
432=>x"0004e",
433=>x"0004e",
434=>x"0004e",
435=>x"0004e",
436=>x"0004e",
437=>x"0004e",
438=>x"0004e",
439=>x"0004e",
440=>x"0004e",
441=>x"0004e",
442=>x"0004e",
443=>x"0004e",
444=>x"0004e",
445=>x"0004e",
446=>x"0004e",
447=>x"0004e",
448=>x"0004e",
449=>x"0004e",
450=>x"0004e",
451=>x"0004e",
452=>x"0004e",
453=>x"0004e",
454=>x"0004f",
455=>x"0004f",
456=>x"0004f",
457=>x"0004f",
458=>x"0004f",
459=>x"0004f",
460=>x"0004f",
461=>x"0004f",
462=>x"0004f",
463=>x"0004f",
464=>x"0004f",
465=>x"0004f",
466=>x"0004f",
467=>x"0004f",
468=>x"0004f",
469=>x"0004f",
470=>x"0004f",
471=>x"0004f",
472=>x"0004f",
473=>x"0004f",
474=>x"0004f",
475=>x"0004f",
476=>x"0004f",
477=>x"0004f",
478=>x"0004f",
479=>x"0004f",
480=>x"0004f",
481=>x"0004f",
482=>x"00050",
483=>x"00050",
484=>x"00050",
485=>x"00050",
486=>x"00050",
487=>x"00050",
488=>x"00050",
489=>x"00050",
490=>x"00050",
491=>x"00050",
492=>x"00050",
493=>x"00050",
494=>x"00050",
495=>x"00050",
496=>x"00050",
497=>x"00050",
498=>x"00050",
499=>x"00050",
500=>x"00050",
501=>x"00050",
502=>x"00050",
503=>x"00050",
504=>x"00050",
505=>x"00050",
506=>x"00050",
507=>x"00050",
508=>x"00050",
509=>x"00050",
510=>x"00050",
511=>x"00050",
512=>x"00051",
513=>x"00051",
514=>x"00051",
515=>x"00051",
516=>x"00051",
517=>x"00051",
518=>x"00051",
519=>x"00051",
520=>x"00051",
521=>x"00051",
522=>x"00051",
523=>x"00051",
524=>x"00051",
525=>x"00051",
526=>x"00051",
527=>x"00051",
528=>x"00051",
529=>x"00051",
530=>x"00051",
531=>x"00051",
532=>x"00051",
533=>x"00051",
534=>x"00051",
535=>x"00051",
536=>x"00051",
537=>x"00051",
538=>x"00051",
539=>x"00051",
540=>x"00051",
541=>x"00051",
542=>x"00051",
543=>x"00051",
544=>x"00051",
545=>x"00051",
546=>x"00052",
547=>x"00052",
548=>x"00052",
549=>x"00052",
550=>x"00052",
551=>x"00052",
552=>x"00052",
553=>x"00052",
554=>x"00052",
555=>x"00052",
556=>x"00052",
557=>x"00052",
558=>x"00052",
559=>x"00052",
560=>x"00052",
561=>x"00052",
562=>x"00052",
563=>x"00052",
564=>x"00052",
565=>x"00052",
566=>x"00052",
567=>x"00052",
568=>x"00052",
569=>x"00052",
570=>x"00052",
571=>x"00052",
572=>x"00052",
573=>x"00052",
574=>x"00052",
575=>x"00052",
576=>x"00052",
577=>x"00052",
578=>x"00052",
579=>x"00052",
580=>x"00052",
581=>x"00052",
582=>x"00052",
583=>x"00052",
584=>x"00053",
585=>x"00053",
586=>x"00053",
587=>x"00053",
588=>x"00053",
589=>x"00053",
590=>x"00053",
591=>x"00053",
592=>x"00053",
593=>x"00053",
594=>x"00053",
595=>x"00053",
596=>x"00053",
597=>x"00053",
598=>x"00053",
599=>x"00053",
600=>x"00053",
601=>x"00053",
602=>x"00053",
603=>x"00053",
604=>x"00053",
605=>x"00053",
606=>x"00053",
607=>x"00053",
608=>x"00053",
609=>x"00053",
610=>x"00053",
611=>x"00053",
612=>x"00053",
613=>x"00053",
614=>x"00053",
615=>x"00053",
616=>x"00053",
617=>x"00053",
618=>x"00053",
619=>x"00053",
620=>x"00053",
621=>x"00053",
622=>x"00053",
623=>x"00053",
624=>x"00053",
625=>x"00054",
626=>x"00054",
627=>x"00054",
628=>x"00054",
629=>x"00054",
630=>x"00054",
631=>x"00054",
632=>x"00054",
633=>x"00054",
634=>x"00054",
635=>x"00054",
636=>x"00054",
637=>x"00054",
638=>x"00054",
639=>x"00054",
640=>x"00054",
641=>x"00054",
642=>x"00054",
643=>x"00054",
644=>x"00054",
645=>x"00054",
646=>x"00054",
647=>x"00054",
648=>x"00054",
649=>x"00054",
650=>x"00054",
651=>x"00054",
652=>x"00054",
653=>x"00054",
654=>x"00054",
655=>x"00054",
656=>x"00054",
657=>x"00054",
658=>x"00054",
659=>x"00054",
660=>x"00054",
661=>x"00054",
662=>x"00054",
663=>x"00054",
664=>x"00054",
665=>x"00054",
666=>x"00054",
667=>x"00054",
668=>x"00054",
669=>x"00054",
670=>x"00054",
671=>x"00054",
672=>x"00055",
673=>x"00055",
674=>x"00055",
675=>x"00055",
676=>x"00055",
677=>x"00055",
678=>x"00055",
679=>x"00055",
680=>x"00055",
681=>x"00055",
682=>x"00055",
683=>x"00055",
684=>x"00055",
685=>x"00055",
686=>x"00055",
687=>x"00055",
688=>x"00055",
689=>x"00055",
690=>x"00055",
691=>x"00055",
692=>x"00055",
693=>x"00055",
694=>x"00055",
695=>x"00055",
696=>x"00055",
697=>x"00055",
698=>x"00055",
699=>x"00055",
700=>x"00055",
701=>x"00055",
702=>x"00055",
703=>x"00055",
704=>x"00055",
705=>x"00055",
706=>x"00055",
707=>x"00055",
708=>x"00055",
709=>x"00055",
710=>x"00055",
711=>x"00055",
712=>x"00055",
713=>x"00055",
714=>x"00055",
715=>x"00055",
716=>x"00055",
717=>x"00055",
718=>x"00055",
719=>x"00055",
720=>x"00055",
721=>x"00055",
722=>x"00055",
723=>x"00055",
724=>x"00055",
725=>x"00055",
726=>x"00056",
727=>x"00056",
728=>x"00056",
729=>x"00056",
730=>x"00056",
731=>x"00056",
732=>x"00056",
733=>x"00056",
734=>x"00056",
735=>x"00056",
736=>x"00056",
737=>x"00056",
738=>x"00056",
739=>x"00056",
740=>x"00056",
741=>x"00056",
742=>x"00056",
743=>x"00056",
744=>x"00056",
745=>x"00056",
746=>x"00056",
747=>x"00056",
748=>x"00056",
749=>x"00056",
750=>x"00056",
751=>x"00056",
752=>x"00056",
753=>x"00056",
754=>x"00056",
755=>x"00056",
756=>x"00056",
757=>x"00056",
758=>x"00056",
759=>x"00056",
760=>x"00056",
761=>x"00056",
762=>x"00056",
763=>x"00056",
764=>x"00056",
765=>x"00056",
766=>x"00056",
767=>x"00056",
768=>x"00056",
769=>x"00056",
770=>x"00056",
771=>x"00056",
772=>x"00056",
773=>x"00056",
774=>x"00056",
775=>x"00056",
776=>x"00056",
777=>x"00056",
778=>x"00056",
779=>x"00056",
780=>x"00056",
781=>x"00056",
782=>x"00056",
783=>x"00056",
784=>x"00056",
785=>x"00056",
786=>x"00056",
787=>x"00057",
788=>x"00057",
789=>x"00057",
790=>x"00057",
791=>x"00057",
792=>x"00057",
793=>x"00057",
794=>x"00057",
795=>x"00057",
796=>x"00057",
797=>x"00057",
798=>x"00057",
799=>x"00057",
800=>x"00057",
801=>x"00057",
802=>x"00057",
803=>x"00057",
804=>x"00057",
805=>x"00057",
806=>x"00057",
807=>x"00057",
808=>x"00057",
809=>x"00057",
810=>x"00057",
811=>x"00057",
812=>x"00057",
813=>x"00057",
814=>x"00057",
815=>x"00057",
816=>x"00057",
817=>x"00057",
818=>x"00057",
819=>x"00057",
820=>x"00057",
821=>x"00057",
822=>x"00057",
823=>x"00057",
824=>x"00057",
825=>x"00057",
826=>x"00057",
827=>x"00057",
828=>x"00057",
829=>x"00057",
830=>x"00057",
831=>x"00057",
832=>x"00057",
833=>x"00057",
834=>x"00057",
835=>x"00057",
836=>x"00057",
837=>x"00057",
838=>x"00057",
839=>x"00057",
840=>x"00057",
841=>x"00057",
842=>x"00057",
843=>x"00057",
844=>x"00057",
845=>x"00057",
846=>x"00057",
847=>x"00057",
848=>x"00057",
849=>x"00057",
850=>x"00057",
851=>x"00057",
852=>x"00057",
853=>x"00057",
854=>x"00057",
855=>x"00057",
856=>x"00057",
857=>x"00058",
858=>x"00058",
859=>x"00058",
860=>x"00058",
861=>x"00058",
862=>x"00058",
863=>x"00058",
864=>x"00058",
865=>x"00058",
866=>x"00058",
867=>x"00058",
868=>x"00058",
869=>x"00058",
870=>x"00058",
871=>x"00058",
872=>x"00058",
873=>x"00058",
874=>x"00058",
875=>x"00058",
876=>x"00058",
877=>x"00058",
878=>x"00058",
879=>x"00058",
880=>x"00058",
881=>x"00058",
882=>x"00058",
883=>x"00058",
884=>x"00058",
885=>x"00058",
886=>x"00058",
887=>x"00058",
888=>x"00058",
889=>x"00058",
890=>x"00058",
891=>x"00058",
892=>x"00058",
893=>x"00058",
894=>x"00058",
895=>x"00058",
896=>x"00058",
897=>x"00058",
898=>x"00058",
899=>x"00058",
900=>x"00058",
901=>x"00058",
902=>x"00058",
903=>x"00058",
904=>x"00058",
905=>x"00058",
906=>x"00058",
907=>x"00058",
908=>x"00058",
909=>x"00058",
910=>x"00058",
911=>x"00058",
912=>x"00058",
913=>x"00058",
914=>x"00058",
915=>x"00058",
916=>x"00058",
917=>x"00058",
918=>x"00058",
919=>x"00058",
920=>x"00058",
921=>x"00058",
922=>x"00058",
923=>x"00058",
924=>x"00058",
925=>x"00058",
926=>x"00058",
927=>x"00058",
928=>x"00058",
929=>x"00058",
930=>x"00058",
931=>x"00058",
932=>x"00058",
933=>x"00058",
934=>x"00058",
935=>x"00058",
936=>x"00058",
937=>x"00058",
938=>x"00058",
939=>x"00059",
940=>x"00059",
941=>x"00059",
942=>x"00059",
943=>x"00059",
944=>x"00059",
945=>x"00059",
946=>x"00059",
947=>x"00059",
948=>x"00059",
949=>x"00059",
950=>x"00059",
951=>x"00059",
952=>x"00059",
953=>x"00059",
954=>x"00059",
955=>x"00059",
956=>x"00059",
957=>x"00059",
958=>x"00059",
959=>x"00059",
960=>x"00059",
961=>x"00059",
962=>x"00059",
963=>x"00059",
964=>x"00059",
965=>x"00059",
966=>x"00059",
967=>x"00059",
968=>x"00059",
969=>x"00059",
970=>x"00059",
971=>x"00059",
972=>x"00059",
973=>x"00059",
974=>x"00059",
975=>x"00059",
976=>x"00059",
977=>x"00059",
978=>x"00059",
979=>x"00059",
980=>x"00059",
981=>x"00059",
982=>x"00059",
983=>x"00059",
984=>x"00059",
985=>x"00059",
986=>x"00059",
987=>x"00059",
988=>x"00059",
989=>x"00059",
990=>x"00059",
991=>x"00059",
992=>x"00059",
993=>x"00059",
994=>x"00059",
995=>x"00059",
996=>x"00059",
997=>x"00059",
998=>x"00059",
999=>x"00059",
1000=>x"00059",
1001=>x"00059",
1002=>x"00059",
1003=>x"00059",
1004=>x"00059",
1005=>x"00059",
1006=>x"00059",
1007=>x"00059",
1008=>x"00059",
1009=>x"00059",
1010=>x"00059",
1011=>x"00059",
1012=>x"00059",
1013=>x"00059",
1014=>x"00059",
1015=>x"00059",
1016=>x"00059",
1017=>x"00059",
1018=>x"00059",
1019=>x"00059",
1020=>x"00059",
1021=>x"00059",
1022=>x"00059",
1023=>x"00059",
1024=>x"00059",
1025=>x"00059",
1026=>x"00059",
1027=>x"00059",
1028=>x"00059",
1029=>x"00059",
1030=>x"00059",
1031=>x"00059",
1032=>x"00059",
1033=>x"00059",
1034=>x"00059",
1035=>x"00059",
1036=>x"0005a",
1037=>x"0005a",
1038=>x"0005a",
1039=>x"0005a",
1040=>x"0005a",
1041=>x"0005a",
1042=>x"0005a",
1043=>x"0005a",
1044=>x"0005a",
1045=>x"0005a",
1046=>x"0005a",
1047=>x"0005a",
1048=>x"0005a",
1049=>x"0005a",
1050=>x"0005a",
1051=>x"0005a",
1052=>x"0005a",
1053=>x"0005a",
1054=>x"0005a",
1055=>x"0005a",
1056=>x"0005a",
1057=>x"0005a",
1058=>x"0005a",
1059=>x"0005a",
1060=>x"0005a",
1061=>x"0005a",
1062=>x"0005a",
1063=>x"0005a",
1064=>x"0005a",
1065=>x"0005a",
1066=>x"0005a",
1067=>x"0005a",
1068=>x"0005a",
1069=>x"0005a",
1070=>x"0005a",
1071=>x"0005a",
1072=>x"0005a",
1073=>x"0005a",
1074=>x"0005a",
1075=>x"0005a",
1076=>x"0005a",
1077=>x"0005a",
1078=>x"0005a",
1079=>x"0005a",
1080=>x"0005a",
1081=>x"0005a",
1082=>x"0005a",
1083=>x"0005a",
1084=>x"0005a",
1085=>x"0005a",
1086=>x"0005a",
1087=>x"0005a",
1088=>x"0005a",
1089=>x"0005a",
1090=>x"0005a",
1091=>x"0005a",
1092=>x"0005a",
1093=>x"0005a",
1094=>x"0005a",
1095=>x"0005a",
1096=>x"0005a",
1097=>x"0005a",
1098=>x"0005a",
1099=>x"0005a",
1100=>x"0005a",
1101=>x"0005a",
1102=>x"0005a",
1103=>x"0005a",
1104=>x"0005a",
1105=>x"0005a",
1106=>x"0005a",
1107=>x"0005a",
1108=>x"0005a",
1109=>x"0005a",
1110=>x"0005a",
1111=>x"0005a",
1112=>x"0005a",
1113=>x"0005a",
1114=>x"0005a",
1115=>x"0005a",
1116=>x"0005a",
1117=>x"0005a",
1118=>x"0005a",
1119=>x"0005a",
1120=>x"0005a",
1121=>x"0005a",
1122=>x"0005a",
1123=>x"0005a",
1124=>x"0005a",
1125=>x"0005a",
1126=>x"0005a",
1127=>x"0005a",
1128=>x"0005a",
1129=>x"0005a",
1130=>x"0005a",
1131=>x"0005a",
1132=>x"0005a",
1133=>x"0005a",
1134=>x"0005a",
1135=>x"0005a",
1136=>x"0005a",
1137=>x"0005a",
1138=>x"0005a",
1139=>x"0005a",
1140=>x"0005a",
1141=>x"0005a",
1142=>x"0005a",
1143=>x"0005a",
1144=>x"0005a",
1145=>x"0005a",
1146=>x"0005a",
1147=>x"0005a",
1148=>x"0005a",
1149=>x"0005a",
1150=>x"0005a",
1151=>x"0005a",
1152=>x"0005b",
1153=>x"0005b",
1154=>x"0005b",
1155=>x"0005b",
1156=>x"0005b",
1157=>x"0005b",
1158=>x"0005b",
1159=>x"0005b",
1160=>x"0005b",
1161=>x"0005b",
1162=>x"0005b",
1163=>x"0005b",
1164=>x"0005b",
1165=>x"0005b",
1166=>x"0005b",
1167=>x"0005b",
1168=>x"0005b",
1169=>x"0005b",
1170=>x"0005b",
1171=>x"0005b",
1172=>x"0005b",
1173=>x"0005b",
1174=>x"0005b",
1175=>x"0005b",
1176=>x"0005b",
1177=>x"0005b",
1178=>x"0005b",
1179=>x"0005b",
1180=>x"0005b",
1181=>x"0005b",
1182=>x"0005b",
1183=>x"0005b",
1184=>x"0005b",
1185=>x"0005b",
1186=>x"0005b",
1187=>x"0005b",
1188=>x"0005b",
1189=>x"0005b",
1190=>x"0005b",
1191=>x"0005b",
1192=>x"0005b",
1193=>x"0005b",
1194=>x"0005b",
1195=>x"0005b",
1196=>x"0005b",
1197=>x"0005b",
1198=>x"0005b",
1199=>x"0005b",
1200=>x"0005b",
1201=>x"0005b",
1202=>x"0005b",
1203=>x"0005b",
1204=>x"0005b",
1205=>x"0005b",
1206=>x"0005b",
1207=>x"0005b",
1208=>x"0005b",
1209=>x"0005b",
1210=>x"0005b",
1211=>x"0005b",
1212=>x"0005b",
1213=>x"0005b",
1214=>x"0005b",
1215=>x"0005b",
1216=>x"0005b",
1217=>x"0005b",
1218=>x"0005b",
1219=>x"0005b",
1220=>x"0005b",
1221=>x"0005b",
1222=>x"0005b",
1223=>x"0005b",
1224=>x"0005b",
1225=>x"0005b",
1226=>x"0005b",
1227=>x"0005b",
1228=>x"0005b",
1229=>x"0005b",
1230=>x"0005b",
1231=>x"0005b",
1232=>x"0005b",
1233=>x"0005b",
1234=>x"0005b",
1235=>x"0005b",
1236=>x"0005b",
1237=>x"0005b",
1238=>x"0005b",
1239=>x"0005b",
1240=>x"0005b",
1241=>x"0005b",
1242=>x"0005b",
1243=>x"0005b",
1244=>x"0005b",
1245=>x"0005b",
1246=>x"0005b",
1247=>x"0005b",
1248=>x"0005b",
1249=>x"0005b",
1250=>x"0005b",
1251=>x"0005b",
1252=>x"0005b",
1253=>x"0005b",
1254=>x"0005b",
1255=>x"0005b",
1256=>x"0005b",
1257=>x"0005b",
1258=>x"0005b",
1259=>x"0005b",
1260=>x"0005b",
1261=>x"0005b",
1262=>x"0005b",
1263=>x"0005b",
1264=>x"0005b",
1265=>x"0005b",
1266=>x"0005b",
1267=>x"0005b",
1268=>x"0005b",
1269=>x"0005b",
1270=>x"0005b",
1271=>x"0005b",
1272=>x"0005b",
1273=>x"0005b",
1274=>x"0005b",
1275=>x"0005b",
1276=>x"0005b",
1277=>x"0005b",
1278=>x"0005b",
1279=>x"0005b",
1280=>x"0005b",
1281=>x"0005b",
1282=>x"0005b",
1283=>x"0005b",
1284=>x"0005b",
1285=>x"0005b",
1286=>x"0005b",
1287=>x"0005b",
1288=>x"0005b",
1289=>x"0005b",
1290=>x"0005b",
1291=>x"0005b",
1292=>x"0005b",
1293=>x"0005b",
1294=>x"0005b",
1295=>x"0005c",
1296=>x"0005c",
1297=>x"0005c",
1298=>x"0005c",
1299=>x"0005c",
1300=>x"0005c",
1301=>x"0005c",
1302=>x"0005c",
1303=>x"0005c",
1304=>x"0005c",
1305=>x"0005c",
1306=>x"0005c",
1307=>x"0005c",
1308=>x"0005c",
1309=>x"0005c",
1310=>x"0005c",
1311=>x"0005c",
1312=>x"0005c",
1313=>x"0005c",
1314=>x"0005c",
1315=>x"0005c",
1316=>x"0005c",
1317=>x"0005c",
1318=>x"0005c",
1319=>x"0005c",
1320=>x"0005c",
1321=>x"0005c",
1322=>x"0005c",
1323=>x"0005c",
1324=>x"0005c",
1325=>x"0005c",
1326=>x"0005c",
1327=>x"0005c",
1328=>x"0005c",
1329=>x"0005c",
1330=>x"0005c",
1331=>x"0005c",
1332=>x"0005c",
1333=>x"0005c",
1334=>x"0005c",
1335=>x"0005c",
1336=>x"0005c",
1337=>x"0005c",
1338=>x"0005c",
1339=>x"0005c",
1340=>x"0005c",
1341=>x"0005c",
1342=>x"0005c",
1343=>x"0005c",
1344=>x"0005c",
1345=>x"0005c",
1346=>x"0005c",
1347=>x"0005c",
1348=>x"0005c",
1349=>x"0005c",
1350=>x"0005c",
1351=>x"0005c",
1352=>x"0005c",
1353=>x"0005c",
1354=>x"0005c",
1355=>x"0005c",
1356=>x"0005c",
1357=>x"0005c",
1358=>x"0005c",
1359=>x"0005c",
1360=>x"0005c",
1361=>x"0005c",
1362=>x"0005c",
1363=>x"0005c",
1364=>x"0005c",
1365=>x"0005c",
1366=>x"0005c",
1367=>x"0005c",
1368=>x"0005c",
1369=>x"0005c",
1370=>x"0005c",
1371=>x"0005c",
1372=>x"0005c",
1373=>x"0005c",
1374=>x"0005c",
1375=>x"0005c",
1376=>x"0005c",
1377=>x"0005c",
1378=>x"0005c",
1379=>x"0005c",
1380=>x"0005c",
1381=>x"0005c",
1382=>x"0005c",
1383=>x"0005c",
1384=>x"0005c",
1385=>x"0005c",
1386=>x"0005c",
1387=>x"0005c",
1388=>x"0005c",
1389=>x"0005c",
1390=>x"0005c",
1391=>x"0005c",
1392=>x"0005c",
1393=>x"0005c",
1394=>x"0005c",
1395=>x"0005c",
1396=>x"0005c",
1397=>x"0005c",
1398=>x"0005c",
1399=>x"0005c",
1400=>x"0005c",
1401=>x"0005c",
1402=>x"0005c",
1403=>x"0005c",
1404=>x"0005c",
1405=>x"0005c",
1406=>x"0005c",
1407=>x"0005c",
1408=>x"0005c",
1409=>x"0005c",
1410=>x"0005c",
1411=>x"0005c",
1412=>x"0005c",
1413=>x"0005c",
1414=>x"0005c",
1415=>x"0005c",
1416=>x"0005c",
1417=>x"0005c",
1418=>x"0005c",
1419=>x"0005c",
1420=>x"0005c",
1421=>x"0005c",
1422=>x"0005c",
1423=>x"0005c",
1424=>x"0005c",
1425=>x"0005c",
1426=>x"0005c",
1427=>x"0005c",
1428=>x"0005c",
1429=>x"0005c",
1430=>x"0005c",
1431=>x"0005c",
1432=>x"0005c",
1433=>x"0005c",
1434=>x"0005c",
1435=>x"0005c",
1436=>x"0005c",
1437=>x"0005c",
1438=>x"0005c",
1439=>x"0005c",
1440=>x"0005c",
1441=>x"0005c",
1442=>x"0005c",
1443=>x"0005c",
1444=>x"0005c",
1445=>x"0005c",
1446=>x"0005c",
1447=>x"0005c",
1448=>x"0005c",
1449=>x"0005c",
1450=>x"0005c",
1451=>x"0005c",
1452=>x"0005c",
1453=>x"0005c",
1454=>x"0005c",
1455=>x"0005c",
1456=>x"0005c",
1457=>x"0005c",
1458=>x"0005c",
1459=>x"0005c",
1460=>x"0005c",
1461=>x"0005c",
1462=>x"0005c",
1463=>x"0005c",
1464=>x"0005c",
1465=>x"0005c",
1466=>x"0005c",
1467=>x"0005c",
1468=>x"0005c",
1469=>x"0005c",
1470=>x"0005c",
1471=>x"0005c",
1472=>x"0005d",
1473=>x"0005d",
1474=>x"0005d",
1475=>x"0005d",
1476=>x"0005d",
1477=>x"0005d",
1478=>x"0005d",
1479=>x"0005d",
1480=>x"0005d",
1481=>x"0005d",
1482=>x"0005d",
1483=>x"0005d",
1484=>x"0005d",
1485=>x"0005d",
1486=>x"0005d",
1487=>x"0005d",
1488=>x"0005d",
1489=>x"0005d",
1490=>x"0005d",
1491=>x"0005d",
1492=>x"0005d",
1493=>x"0005d",
1494=>x"0005d",
1495=>x"0005d",
1496=>x"0005d",
1497=>x"0005d",
1498=>x"0005d",
1499=>x"0005d",
1500=>x"0005d",
1501=>x"0005d",
1502=>x"0005d",
1503=>x"0005d",
1504=>x"0005d",
1505=>x"0005d",
1506=>x"0005d",
1507=>x"0005d",
1508=>x"0005d",
1509=>x"0005d",
1510=>x"0005d",
1511=>x"0005d",
1512=>x"0005d",
1513=>x"0005d",
1514=>x"0005d",
1515=>x"0005d",
1516=>x"0005d",
1517=>x"0005d",
1518=>x"0005d",
1519=>x"0005d",
1520=>x"0005d",
1521=>x"0005d",
1522=>x"0005d",
1523=>x"0005d",
1524=>x"0005d",
1525=>x"0005d",
1526=>x"0005d",
1527=>x"0005d",
1528=>x"0005d",
1529=>x"0005d",
1530=>x"0005d",
1531=>x"0005d",
1532=>x"0005d",
1533=>x"0005d",
1534=>x"0005d",
1535=>x"0005d",
1536=>x"0005d",
1537=>x"0005d",
1538=>x"0005d",
1539=>x"0005d",
1540=>x"0005d",
1541=>x"0005d",
1542=>x"0005d",
1543=>x"0005d",
1544=>x"0005d",
1545=>x"0005d",
1546=>x"0005d",
1547=>x"0005d",
1548=>x"0005d",
1549=>x"0005d",
1550=>x"0005d",
1551=>x"0005d",
1552=>x"0005d",
1553=>x"0005d",
1554=>x"0005d",
1555=>x"0005d",
1556=>x"0005d",
1557=>x"0005d",
1558=>x"0005d",
1559=>x"0005d",
1560=>x"0005d",
1561=>x"0005d",
1562=>x"0005d",
1563=>x"0005d",
1564=>x"0005d",
1565=>x"0005d",
1566=>x"0005d",
1567=>x"0005d",
1568=>x"0005d",
1569=>x"0005d",
1570=>x"0005d",
1571=>x"0005d",
1572=>x"0005d",
1573=>x"0005d",
1574=>x"0005d",
1575=>x"0005d",
1576=>x"0005d",
1577=>x"0005d",
1578=>x"0005d",
1579=>x"0005d",
1580=>x"0005d",
1581=>x"0005d",
1582=>x"0005d",
1583=>x"0005d",
1584=>x"0005d",
1585=>x"0005d",
1586=>x"0005d",
1587=>x"0005d",
1588=>x"0005d",
1589=>x"0005d",
1590=>x"0005d",
1591=>x"0005d",
1592=>x"0005d",
1593=>x"0005d",
1594=>x"0005d",
1595=>x"0005d",
1596=>x"0005d",
1597=>x"0005d",
1598=>x"0005d",
1599=>x"0005d",
1600=>x"0005d",
1601=>x"0005d",
1602=>x"0005d",
1603=>x"0005d",
1604=>x"0005d",
1605=>x"0005d",
1606=>x"0005d",
1607=>x"0005d",
1608=>x"0005d",
1609=>x"0005d",
1610=>x"0005d",
1611=>x"0005d",
1612=>x"0005d",
1613=>x"0005d",
1614=>x"0005d",
1615=>x"0005d",
1616=>x"0005d",
1617=>x"0005d",
1618=>x"0005d",
1619=>x"0005d",
1620=>x"0005d",
1621=>x"0005d",
1622=>x"0005d",
1623=>x"0005d",
1624=>x"0005d",
1625=>x"0005d",
1626=>x"0005d",
1627=>x"0005d",
1628=>x"0005d",
1629=>x"0005d",
1630=>x"0005d",
1631=>x"0005d",
1632=>x"0005d",
1633=>x"0005d",
1634=>x"0005d",
1635=>x"0005d",
1636=>x"0005d",
1637=>x"0005d",
1638=>x"0005d",
1639=>x"0005d",
1640=>x"0005d",
1641=>x"0005d",
1642=>x"0005d",
1643=>x"0005d",
1644=>x"0005d",
1645=>x"0005d",
1646=>x"0005d",
1647=>x"0005d",
1648=>x"0005d",
1649=>x"0005d",
1650=>x"0005d",
1651=>x"0005d",
1652=>x"0005d",
1653=>x"0005d",
1654=>x"0005d",
1655=>x"0005d",
1656=>x"0005d",
1657=>x"0005d",
1658=>x"0005d",
1659=>x"0005d",
1660=>x"0005d",
1661=>x"0005d",
1662=>x"0005d",
1663=>x"0005d",
1664=>x"0005d",
1665=>x"0005d",
1666=>x"0005d",
1667=>x"0005d",
1668=>x"0005d",
1669=>x"0005d",
1670=>x"0005d",
1671=>x"0005d",
1672=>x"0005d",
1673=>x"0005d",
1674=>x"0005d",
1675=>x"0005d",
1676=>x"0005d",
1677=>x"0005d",
1678=>x"0005d",
1679=>x"0005d",
1680=>x"0005d",
1681=>x"0005d",
1682=>x"0005d",
1683=>x"0005d",
1684=>x"0005d",
1685=>x"0005d",
1686=>x"0005d",
1687=>x"0005d",
1688=>x"0005d",
1689=>x"0005d",
1690=>x"0005d",
1691=>x"0005d",
1692=>x"0005d",
1693=>x"0005d",
1694=>x"0005d",
1695=>x"0005d",
1696=>x"0005d",
1697=>x"0005d",
1698=>x"0005d",
1699=>x"0005d",
1700=>x"0005d",
1701=>x"0005e",
1702=>x"0005e",
1703=>x"0005e",
1704=>x"0005e",
1705=>x"0005e",
1706=>x"0005e",
1707=>x"0005e",
1708=>x"0005e",
1709=>x"0005e",
1710=>x"0005e",
1711=>x"0005e",
1712=>x"0005e",
1713=>x"0005e",
1714=>x"0005e",
1715=>x"0005e",
1716=>x"0005e",
1717=>x"0005e",
1718=>x"0005e",
1719=>x"0005e",
1720=>x"0005e",
1721=>x"0005e",
1722=>x"0005e",
1723=>x"0005e",
1724=>x"0005e",
1725=>x"0005e",
1726=>x"0005e",
1727=>x"0005e",
1728=>x"0005e",
1729=>x"0005e",
1730=>x"0005e",
1731=>x"0005e",
1732=>x"0005e",
1733=>x"0005e",
1734=>x"0005e",
1735=>x"0005e",
1736=>x"0005e",
1737=>x"0005e",
1738=>x"0005e",
1739=>x"0005e",
1740=>x"0005e",
1741=>x"0005e",
1742=>x"0005e",
1743=>x"0005e",
1744=>x"0005e",
1745=>x"0005e",
1746=>x"0005e",
1747=>x"0005e",
1748=>x"0005e",
1749=>x"0005e",
1750=>x"0005e",
1751=>x"0005e",
1752=>x"0005e",
1753=>x"0005e",
1754=>x"0005e",
1755=>x"0005e",
1756=>x"0005e",
1757=>x"0005e",
1758=>x"0005e",
1759=>x"0005e",
1760=>x"0005e",
1761=>x"0005e",
1762=>x"0005e",
1763=>x"0005e",
1764=>x"0005e",
1765=>x"0005e",
1766=>x"0005e",
1767=>x"0005e",
1768=>x"0005e",
1769=>x"0005e",
1770=>x"0005e",
1771=>x"0005e",
1772=>x"0005e",
1773=>x"0005e",
1774=>x"0005e",
1775=>x"0005e",
1776=>x"0005e",
1777=>x"0005e",
1778=>x"0005e",
1779=>x"0005e",
1780=>x"0005e",
1781=>x"0005e",
1782=>x"0005e",
1783=>x"0005e",
1784=>x"0005e",
1785=>x"0005e",
1786=>x"0005e",
1787=>x"0005e",
1788=>x"0005e",
1789=>x"0005e",
1790=>x"0005e",
1791=>x"0005e",
1792=>x"0005e",
1793=>x"0005e",
1794=>x"0005e",
1795=>x"0005e",
1796=>x"0005e",
1797=>x"0005e",
1798=>x"0005e",
1799=>x"0005e",
1800=>x"0005e",
1801=>x"0005e",
1802=>x"0005e",
1803=>x"0005e",
1804=>x"0005e",
1805=>x"0005e",
1806=>x"0005e",
1807=>x"0005e",
1808=>x"0005e",
1809=>x"0005e",
1810=>x"0005e",
1811=>x"0005e",
1812=>x"0005e",
1813=>x"0005e",
1814=>x"0005e",
1815=>x"0005e",
1816=>x"0005e",
1817=>x"0005e",
1818=>x"0005e",
1819=>x"0005e",
1820=>x"0005e",
1821=>x"0005e",
1822=>x"0005e",
1823=>x"0005e",
1824=>x"0005e",
1825=>x"0005e",
1826=>x"0005e",
1827=>x"0005e",
1828=>x"0005e",
1829=>x"0005e",
1830=>x"0005e",
1831=>x"0005e",
1832=>x"0005e",
1833=>x"0005e",
1834=>x"0005e",
1835=>x"0005e",
1836=>x"0005e",
1837=>x"0005e",
1838=>x"0005e",
1839=>x"0005e",
1840=>x"0005e",
1841=>x"0005e",
1842=>x"0005e",
1843=>x"0005e",
1844=>x"0005e",
1845=>x"0005e",
1846=>x"0005e",
1847=>x"0005e",
1848=>x"0005e",
1849=>x"0005e",
1850=>x"0005e",
1851=>x"0005e",
1852=>x"0005e",
1853=>x"0005e",
1854=>x"0005e",
1855=>x"0005e",
1856=>x"0005e",
1857=>x"0005e",
1858=>x"0005e",
1859=>x"0005e",
1860=>x"0005e",
1861=>x"0005e",
1862=>x"0005e",
1863=>x"0005e",
1864=>x"0005e",
1865=>x"0005e",
1866=>x"0005e",
1867=>x"0005e",
1868=>x"0005e",
1869=>x"0005e",
1870=>x"0005e",
1871=>x"0005e",
1872=>x"0005e",
1873=>x"0005e",
1874=>x"0005e",
1875=>x"0005e",
1876=>x"0005e",
1877=>x"0005e",
1878=>x"0005e",
1879=>x"0005e",
1880=>x"0005e",
1881=>x"0005e",
1882=>x"0005e",
1883=>x"0005e",
1884=>x"0005e",
1885=>x"0005e",
1886=>x"0005e",
1887=>x"0005e",
1888=>x"0005e",
1889=>x"0005e",
1890=>x"0005e",
1891=>x"0005e",
1892=>x"0005e",
1893=>x"0005e",
1894=>x"0005e",
1895=>x"0005e",
1896=>x"0005e",
1897=>x"0005e",
1898=>x"0005e",
1899=>x"0005e",
1900=>x"0005e",
1901=>x"0005e",
1902=>x"0005e",
1903=>x"0005e",
1904=>x"0005e",
1905=>x"0005e",
1906=>x"0005e",
1907=>x"0005e",
1908=>x"0005e",
1909=>x"0005e",
1910=>x"0005e",
1911=>x"0005e",
1912=>x"0005e",
1913=>x"0005e",
1914=>x"0005e",
1915=>x"0005e",
1916=>x"0005e",
1917=>x"0005e",
1918=>x"0005e",
1919=>x"0005e",
1920=>x"0005e",
1921=>x"0005e",
1922=>x"0005e",
1923=>x"0005e",
1924=>x"0005e",
1925=>x"0005e",
1926=>x"0005e",
1927=>x"0005e",
1928=>x"0005e",
1929=>x"0005e",
1930=>x"0005e",
1931=>x"0005e",
1932=>x"0005e",
1933=>x"0005e",
1934=>x"0005e",
1935=>x"0005e",
1936=>x"0005e",
1937=>x"0005e",
1938=>x"0005e",
1939=>x"0005e",
1940=>x"0005e",
1941=>x"0005e",
1942=>x"0005e",
1943=>x"0005e",
1944=>x"0005e",
1945=>x"0005e",
1946=>x"0005e",
1947=>x"0005e",
1948=>x"0005e",
1949=>x"0005e",
1950=>x"0005e",
1951=>x"0005e",
1952=>x"0005e",
1953=>x"0005e",
1954=>x"0005e",
1955=>x"0005e",
1956=>x"0005e",
1957=>x"0005e",
1958=>x"0005e",
1959=>x"0005e",
1960=>x"0005e",
1961=>x"0005e",
1962=>x"0005e",
1963=>x"0005e",
1964=>x"0005e",
1965=>x"0005e",
1966=>x"0005e",
1967=>x"0005e",
1968=>x"0005e",
1969=>x"0005e",
1970=>x"0005e",
1971=>x"0005e",
1972=>x"0005e",
1973=>x"0005e",
1974=>x"0005e",
1975=>x"0005e",
1976=>x"0005e",
1977=>x"0005e",
1978=>x"0005e",
1979=>x"0005e",
1980=>x"0005e",
1981=>x"0005e",
1982=>x"0005e",
1983=>x"0005e",
1984=>x"0005e",
1985=>x"0005e",
1986=>x"0005e",
1987=>x"0005e",
1988=>x"0005e",
1989=>x"0005e",
1990=>x"0005e",
1991=>x"0005e",
1992=>x"0005e",
1993=>x"0005e",
1994=>x"0005e",
1995=>x"0005e",
1996=>x"0005e",
1997=>x"0005e",
1998=>x"0005e",
1999=>x"0005e",
2000=>x"0005e",
2001=>x"0005e",
2002=>x"0005e",
2003=>x"0005e",
2004=>x"0005e",
2005=>x"0005e",
2006=>x"0005f",
2007=>x"0005f",
2008=>x"0005f",
2009=>x"0005f",
2010=>x"0005f",
2011=>x"0005f",
2012=>x"0005f",
2013=>x"0005f",
2014=>x"0005f",
2015=>x"0005f",
2016=>x"0005f",
2017=>x"0005f",
2018=>x"0005f",
2019=>x"0005f",
2020=>x"0005f",
2021=>x"0005f",
2022=>x"0005f",
2023=>x"0005f",
2024=>x"0005f",
2025=>x"0005f",
2026=>x"0005f",
2027=>x"0005f",
2028=>x"0005f",
2029=>x"0005f",
2030=>x"0005f",
2031=>x"0005f",
2032=>x"0005f",
2033=>x"0005f",
2034=>x"0005f",
2035=>x"0005f",
2036=>x"0005f",
2037=>x"0005f",
2038=>x"0005f",
2039=>x"0005f",
2040=>x"0005f",
2041=>x"0005f",
2042=>x"0005f",
2043=>x"0005f",
2044=>x"0005f",
2045=>x"0005f",
2046=>x"0005f",
2047=>x"0005f",
2048=>x"0005f",
2049=>x"0005f",
2050=>x"0005f",
2051=>x"0005f",
2052=>x"0005f",
2053=>x"0005f",
2054=>x"0005f",
2055=>x"0005f",
2056=>x"0005f",
2057=>x"0005f",
2058=>x"0005f",
2059=>x"0005f",
2060=>x"0005f",
2061=>x"0005f",
2062=>x"0005f",
2063=>x"0005f",
2064=>x"0005f",
2065=>x"0005f",
2066=>x"0005f",
2067=>x"0005f",
2068=>x"0005f",
2069=>x"0005f",
2070=>x"0005f",
2071=>x"0005f",
2072=>x"0005f",
2073=>x"0005f",
2074=>x"0005f",
2075=>x"0005f",
2076=>x"0005f",
2077=>x"0005f",
2078=>x"0005f",
2079=>x"0005f",
2080=>x"0005f",
2081=>x"0005f",
2082=>x"0005f",
2083=>x"0005f",
2084=>x"0005f",
2085=>x"0005f",
2086=>x"0005f",
2087=>x"0005f",
2088=>x"0005f",
2089=>x"0005f",
2090=>x"0005f",
2091=>x"0005f",
2092=>x"0005f",
2093=>x"0005f",
2094=>x"0005f",
2095=>x"0005f",
2096=>x"0005f",
2097=>x"0005f",
2098=>x"0005f",
2099=>x"0005f",
2100=>x"0005f",
2101=>x"0005f",
2102=>x"0005f",
2103=>x"0005f",
2104=>x"0005f",
2105=>x"0005f",
2106=>x"0005f",
2107=>x"0005f",
2108=>x"0005f",
2109=>x"0005f",
2110=>x"0005f",
2111=>x"0005f",
2112=>x"0005f",
2113=>x"0005f",
2114=>x"0005f",
2115=>x"0005f",
2116=>x"0005f",
2117=>x"0005f",
2118=>x"0005f",
2119=>x"0005f",
2120=>x"0005f",
2121=>x"0005f",
2122=>x"0005f",
2123=>x"0005f",
2124=>x"0005f",
2125=>x"0005f",
2126=>x"0005f",
2127=>x"0005f",
2128=>x"0005f",
2129=>x"0005f",
2130=>x"0005f",
2131=>x"0005f",
2132=>x"0005f",
2133=>x"0005f",
2134=>x"0005f",
2135=>x"0005f",
2136=>x"0005f",
2137=>x"0005f",
2138=>x"0005f",
2139=>x"0005f",
2140=>x"0005f",
2141=>x"0005f",
2142=>x"0005f",
2143=>x"0005f",
2144=>x"0005f",
2145=>x"0005f",
2146=>x"0005f",
2147=>x"0005f",
2148=>x"0005f",
2149=>x"0005f",
2150=>x"0005f",
2151=>x"0005f",
2152=>x"0005f",
2153=>x"0005f",
2154=>x"0005f",
2155=>x"0005f",
2156=>x"0005f",
2157=>x"0005f",
2158=>x"0005f",
2159=>x"0005f",
2160=>x"0005f",
2161=>x"0005f",
2162=>x"0005f",
2163=>x"0005f",
2164=>x"0005f",
2165=>x"0005f",
2166=>x"0005f",
2167=>x"0005f",
2168=>x"0005f",
2169=>x"0005f",
2170=>x"0005f",
2171=>x"0005f",
2172=>x"0005f",
2173=>x"0005f",
2174=>x"0005f",
2175=>x"0005f",
2176=>x"0005f",
2177=>x"0005f",
2178=>x"0005f",
2179=>x"0005f",
2180=>x"0005f",
2181=>x"0005f",
2182=>x"0005f",
2183=>x"0005f",
2184=>x"0005f",
2185=>x"0005f",
2186=>x"0005f",
2187=>x"0005f",
2188=>x"0005f",
2189=>x"0005f",
2190=>x"0005f",
2191=>x"0005f",
2192=>x"0005f",
2193=>x"0005f",
2194=>x"0005f",
2195=>x"0005f",
2196=>x"0005f",
2197=>x"0005f",
2198=>x"0005f",
2199=>x"0005f",
2200=>x"0005f",
2201=>x"0005f",
2202=>x"0005f",
2203=>x"0005f",
2204=>x"0005f",
2205=>x"0005f",
2206=>x"0005f",
2207=>x"0005f",
2208=>x"0005f",
2209=>x"0005f",
2210=>x"0005f",
2211=>x"0005f",
2212=>x"0005f",
2213=>x"0005f",
2214=>x"0005f",
2215=>x"0005f",
2216=>x"0005f",
2217=>x"0005f",
2218=>x"0005f",
2219=>x"0005f",
2220=>x"0005f",
2221=>x"0005f",
2222=>x"0005f",
2223=>x"0005f",
2224=>x"0005f",
2225=>x"0005f",
2226=>x"0005f",
2227=>x"0005f",
2228=>x"0005f",
2229=>x"0005f",
2230=>x"0005f",
2231=>x"0005f",
2232=>x"0005f",
2233=>x"0005f",
2234=>x"0005f",
2235=>x"0005f",
2236=>x"0005f",
2237=>x"0005f",
2238=>x"0005f",
2239=>x"0005f",
2240=>x"0005f",
2241=>x"0005f",
2242=>x"0005f",
2243=>x"0005f",
2244=>x"0005f",
2245=>x"0005f",
2246=>x"0005f",
2247=>x"0005f",
2248=>x"0005f",
2249=>x"0005f",
2250=>x"0005f",
2251=>x"0005f",
2252=>x"0005f",
2253=>x"0005f",
2254=>x"0005f",
2255=>x"0005f",
2256=>x"0005f",
2257=>x"0005f",
2258=>x"0005f",
2259=>x"0005f",
2260=>x"0005f",
2261=>x"0005f",
2262=>x"0005f",
2263=>x"0005f",
2264=>x"0005f",
2265=>x"0005f",
2266=>x"0005f",
2267=>x"0005f",
2268=>x"0005f",
2269=>x"0005f",
2270=>x"0005f",
2271=>x"0005f",
2272=>x"0005f",
2273=>x"0005f",
2274=>x"0005f",
2275=>x"0005f",
2276=>x"0005f",
2277=>x"0005f",
2278=>x"0005f",
2279=>x"0005f",
2280=>x"0005f",
2281=>x"0005f",
2282=>x"0005f",
2283=>x"0005f",
2284=>x"0005f",
2285=>x"0005f",
2286=>x"0005f",
2287=>x"0005f",
2288=>x"0005f",
2289=>x"0005f",
2290=>x"0005f",
2291=>x"0005f",
2292=>x"0005f",
2293=>x"0005f",
2294=>x"0005f",
2295=>x"0005f",
2296=>x"0005f",
2297=>x"0005f",
2298=>x"0005f",
2299=>x"0005f",
2300=>x"0005f",
2301=>x"0005f",
2302=>x"0005f",
2303=>x"0005f",
2304=>x"0005f",
2305=>x"0005f",
2306=>x"0005f",
2307=>x"0005f",
2308=>x"0005f",
2309=>x"0005f",
2310=>x"0005f",
2311=>x"0005f",
2312=>x"0005f",
2313=>x"0005f",
2314=>x"0005f",
2315=>x"0005f",
2316=>x"0005f",
2317=>x"0005f",
2318=>x"0005f",
2319=>x"0005f",
2320=>x"0005f",
2321=>x"0005f",
2322=>x"0005f",
2323=>x"0005f",
2324=>x"0005f",
2325=>x"0005f",
2326=>x"0005f",
2327=>x"0005f",
2328=>x"0005f",
2329=>x"0005f",
2330=>x"0005f",
2331=>x"0005f",
2332=>x"0005f",
2333=>x"0005f",
2334=>x"0005f",
2335=>x"0005f",
2336=>x"0005f",
2337=>x"0005f",
2338=>x"0005f",
2339=>x"0005f",
2340=>x"0005f",
2341=>x"0005f",
2342=>x"0005f",
2343=>x"0005f",
2344=>x"0005f",
2345=>x"0005f",
2346=>x"0005f",
2347=>x"0005f",
2348=>x"0005f",
2349=>x"0005f",
2350=>x"0005f",
2351=>x"0005f",
2352=>x"0005f",
2353=>x"0005f",
2354=>x"0005f",
2355=>x"0005f",
2356=>x"0005f",
2357=>x"0005f",
2358=>x"0005f",
2359=>x"0005f",
2360=>x"0005f",
2361=>x"0005f",
2362=>x"0005f",
2363=>x"0005f",
2364=>x"0005f",
2365=>x"0005f",
2366=>x"0005f",
2367=>x"0005f",
2368=>x"0005f",
2369=>x"0005f",
2370=>x"0005f",
2371=>x"0005f",
2372=>x"0005f",
2373=>x"0005f",
2374=>x"0005f",
2375=>x"0005f",
2376=>x"0005f",
2377=>x"0005f",
2378=>x"0005f",
2379=>x"0005f",
2380=>x"0005f",
2381=>x"0005f",
2382=>x"0005f",
2383=>x"0005f",
2384=>x"0005f",
2385=>x"0005f",
2386=>x"0005f",
2387=>x"0005f",
2388=>x"0005f",
2389=>x"0005f",
2390=>x"0005f",
2391=>x"0005f",
2392=>x"0005f",
2393=>x"0005f",
2394=>x"0005f",
2395=>x"0005f",
2396=>x"0005f",
2397=>x"0005f",
2398=>x"0005f",
2399=>x"0005f",
2400=>x"0005f",
2401=>x"0005f",
2402=>x"0005f",
2403=>x"0005f",
2404=>x"0005f",
2405=>x"0005f",
2406=>x"0005f",
2407=>x"0005f",
2408=>x"0005f",
2409=>x"0005f",
2410=>x"0005f",
2411=>x"0005f",
2412=>x"0005f",
2413=>x"0005f",
2414=>x"0005f",
2415=>x"0005f",
2416=>x"0005f",
2417=>x"0005f",
2418=>x"0005f",
2419=>x"0005f",
2420=>x"0005f",
2421=>x"0005f",
2422=>x"0005f",
2423=>x"0005f",
2424=>x"0005f",
2425=>x"0005f",
2426=>x"0005f",
2427=>x"0005f",
2428=>x"0005f",
2429=>x"0005f",
2430=>x"0005f",
2431=>x"0005f",
2432=>x"00060",
2433=>x"00060",
2434=>x"00060",
2435=>x"00060",
2436=>x"00060",
2437=>x"00060",
2438=>x"00060",
2439=>x"00060",
2440=>x"00060",
2441=>x"00060",
2442=>x"00060",
2443=>x"00060",
2444=>x"00060",
2445=>x"00060",
2446=>x"00060",
2447=>x"00060",
2448=>x"00060",
2449=>x"00060",
2450=>x"00060",
2451=>x"00060",
2452=>x"00060",
2453=>x"00060",
2454=>x"00060",
2455=>x"00060",
2456=>x"00060",
2457=>x"00060",
2458=>x"00060",
2459=>x"00060",
2460=>x"00060",
2461=>x"00060",
2462=>x"00060",
2463=>x"00060",
2464=>x"00060",
2465=>x"00060",
2466=>x"00060",
2467=>x"00060",
2468=>x"00060",
2469=>x"00060",
2470=>x"00060",
2471=>x"00060",
2472=>x"00060",
2473=>x"00060",
2474=>x"00060",
2475=>x"00060",
2476=>x"00060",
2477=>x"00060",
2478=>x"00060",
2479=>x"00060",
2480=>x"00060",
2481=>x"00060",
2482=>x"00060",
2483=>x"00060",
2484=>x"00060",
2485=>x"00060",
2486=>x"00060",
2487=>x"00060",
2488=>x"00060",
2489=>x"00060",
2490=>x"00060",
2491=>x"00060",
2492=>x"00060",
2493=>x"00060",
2494=>x"00060",
2495=>x"00060",
2496=>x"00060",
2497=>x"00060",
2498=>x"00060",
2499=>x"00060",
2500=>x"00060",
2501=>x"00060",
2502=>x"00060",
2503=>x"00060",
2504=>x"00060",
2505=>x"00060",
2506=>x"00060",
2507=>x"00060",
2508=>x"00060",
2509=>x"00060",
2510=>x"00060",
2511=>x"00060",
2512=>x"00060",
2513=>x"00060",
2514=>x"00060",
2515=>x"00060",
2516=>x"00060",
2517=>x"00060",
2518=>x"00060",
2519=>x"00060",
2520=>x"00060",
2521=>x"00060",
2522=>x"00060",
2523=>x"00060",
2524=>x"00060",
2525=>x"00060",
2526=>x"00060",
2527=>x"00060",
2528=>x"00060",
2529=>x"00060",
2530=>x"00060",
2531=>x"00060",
2532=>x"00060",
2533=>x"00060",
2534=>x"00060",
2535=>x"00060",
2536=>x"00060",
2537=>x"00060",
2538=>x"00060",
2539=>x"00060",
2540=>x"00060",
2541=>x"00060",
2542=>x"00060",
2543=>x"00060",
2544=>x"00060",
2545=>x"00060",
2546=>x"00060",
2547=>x"00060",
2548=>x"00060",
2549=>x"00060",
2550=>x"00060",
2551=>x"00060",
2552=>x"00060",
2553=>x"00060",
2554=>x"00060",
2555=>x"00060",
2556=>x"00060",
2557=>x"00060",
2558=>x"00060",
2559=>x"00060",
2560=>x"00060",
2561=>x"00060",
2562=>x"00060",
2563=>x"00060",
2564=>x"00060",
2565=>x"00060",
2566=>x"00060",
2567=>x"00060",
2568=>x"00060",
2569=>x"00060",
2570=>x"00060",
2571=>x"00060",
2572=>x"00060",
2573=>x"00060",
2574=>x"00060",
2575=>x"00060",
2576=>x"00060",
2577=>x"00060",
2578=>x"00060",
2579=>x"00060",
2580=>x"00060",
2581=>x"00060",
2582=>x"00060",
2583=>x"00060",
2584=>x"00060",
2585=>x"00060",
2586=>x"00060",
2587=>x"00060",
2588=>x"00060",
2589=>x"00060",
2590=>x"00060",
2591=>x"00060",
2592=>x"00060",
2593=>x"00060",
2594=>x"00060",
2595=>x"00060",
2596=>x"00060",
2597=>x"00060",
2598=>x"00060",
2599=>x"00060",
2600=>x"00060",
2601=>x"00060",
2602=>x"00060",
2603=>x"00060",
2604=>x"00060",
2605=>x"00060",
2606=>x"00060",
2607=>x"00060",
2608=>x"00060",
2609=>x"00060",
2610=>x"00060",
2611=>x"00060",
2612=>x"00060",
2613=>x"00060",
2614=>x"00060",
2615=>x"00060",
2616=>x"00060",
2617=>x"00060",
2618=>x"00060",
2619=>x"00060",
2620=>x"00060",
2621=>x"00060",
2622=>x"00060",
2623=>x"00060",
2624=>x"00060",
2625=>x"00060",
2626=>x"00060",
2627=>x"00060",
2628=>x"00060",
2629=>x"00060",
2630=>x"00060",
2631=>x"00060",
2632=>x"00060",
2633=>x"00060",
2634=>x"00060",
2635=>x"00060",
2636=>x"00060",
2637=>x"00060",
2638=>x"00060",
2639=>x"00060",
2640=>x"00060",
2641=>x"00060",
2642=>x"00060",
2643=>x"00060",
2644=>x"00060",
2645=>x"00060",
2646=>x"00060",
2647=>x"00060",
2648=>x"00060",
2649=>x"00060",
2650=>x"00060",
2651=>x"00060",
2652=>x"00060",
2653=>x"00060",
2654=>x"00060",
2655=>x"00060",
2656=>x"00060",
2657=>x"00060",
2658=>x"00060",
2659=>x"00060",
2660=>x"00060",
2661=>x"00060",
2662=>x"00060",
2663=>x"00060",
2664=>x"00060",
2665=>x"00060",
2666=>x"00060",
2667=>x"00060",
2668=>x"00060",
2669=>x"00060",
2670=>x"00060",
2671=>x"00060",
2672=>x"00060",
2673=>x"00060",
2674=>x"00060",
2675=>x"00060",
2676=>x"00060",
2677=>x"00060",
2678=>x"00060",
2679=>x"00060",
2680=>x"00060",
2681=>x"00060",
2682=>x"00060",
2683=>x"00060",
2684=>x"00060",
2685=>x"00060",
2686=>x"00060",
2687=>x"00060",
2688=>x"00060",
2689=>x"00060",
2690=>x"00060",
2691=>x"00060",
2692=>x"00060",
2693=>x"00060",
2694=>x"00060",
2695=>x"00060",
2696=>x"00060",
2697=>x"00060",
2698=>x"00060",
2699=>x"00060",
2700=>x"00060",
2701=>x"00060",
2702=>x"00060",
2703=>x"00060",
2704=>x"00060",
2705=>x"00060",
2706=>x"00060",
2707=>x"00060",
2708=>x"00060",
2709=>x"00060",
2710=>x"00060",
2711=>x"00060",
2712=>x"00060",
2713=>x"00060",
2714=>x"00060",
2715=>x"00060",
2716=>x"00060",
2717=>x"00060",
2718=>x"00060",
2719=>x"00060",
2720=>x"00060",
2721=>x"00060",
2722=>x"00060",
2723=>x"00060",
2724=>x"00060",
2725=>x"00060",
2726=>x"00060",
2727=>x"00060",
2728=>x"00060",
2729=>x"00060",
2730=>x"00060",
2731=>x"00060",
2732=>x"00060",
2733=>x"00060",
2734=>x"00060",
2735=>x"00060",
2736=>x"00060",
2737=>x"00060",
2738=>x"00060",
2739=>x"00060",
2740=>x"00060",
2741=>x"00060",
2742=>x"00060",
2743=>x"00060",
2744=>x"00060",
2745=>x"00060",
2746=>x"00060",
2747=>x"00060",
2748=>x"00060",
2749=>x"00060",
2750=>x"00060",
2751=>x"00060",
2752=>x"00060",
2753=>x"00060",
2754=>x"00060",
2755=>x"00060",
2756=>x"00060",
2757=>x"00060",
2758=>x"00060",
2759=>x"00060",
2760=>x"00060",
2761=>x"00060",
2762=>x"00060",
2763=>x"00060",
2764=>x"00060",
2765=>x"00060",
2766=>x"00060",
2767=>x"00060",
2768=>x"00060",
2769=>x"00060",
2770=>x"00060",
2771=>x"00060",
2772=>x"00060",
2773=>x"00060",
2774=>x"00060",
2775=>x"00060",
2776=>x"00060",
2777=>x"00060",
2778=>x"00060",
2779=>x"00060",
2780=>x"00060",
2781=>x"00060",
2782=>x"00060",
2783=>x"00060",
2784=>x"00060",
2785=>x"00060",
2786=>x"00060",
2787=>x"00060",
2788=>x"00060",
2789=>x"00060",
2790=>x"00060",
2791=>x"00060",
2792=>x"00060",
2793=>x"00060",
2794=>x"00060",
2795=>x"00060",
2796=>x"00060",
2797=>x"00060",
2798=>x"00060",
2799=>x"00060",
2800=>x"00060",
2801=>x"00060",
2802=>x"00060",
2803=>x"00060",
2804=>x"00060",
2805=>x"00060",
2806=>x"00060",
2807=>x"00060",
2808=>x"00060",
2809=>x"00060",
2810=>x"00060",
2811=>x"00060",
2812=>x"00060",
2813=>x"00060",
2814=>x"00060",
2815=>x"00060",
2816=>x"00060",
2817=>x"00060",
2818=>x"00060",
2819=>x"00060",
2820=>x"00060",
2821=>x"00060",
2822=>x"00060",
2823=>x"00060",
2824=>x"00060",
2825=>x"00060",
2826=>x"00060",
2827=>x"00060",
2828=>x"00060",
2829=>x"00060",
2830=>x"00060",
2831=>x"00060",
2832=>x"00060",
2833=>x"00060",
2834=>x"00060",
2835=>x"00060",
2836=>x"00060",
2837=>x"00060",
2838=>x"00060",
2839=>x"00060",
2840=>x"00060",
2841=>x"00060",
2842=>x"00060",
2843=>x"00060",
2844=>x"00060",
2845=>x"00060",
2846=>x"00060",
2847=>x"00060",
2848=>x"00060",
2849=>x"00060",
2850=>x"00060",
2851=>x"00060",
2852=>x"00060",
2853=>x"00060",
2854=>x"00060",
2855=>x"00060",
2856=>x"00060",
2857=>x"00060",
2858=>x"00060",
2859=>x"00060",
2860=>x"00060",
2861=>x"00060",
2862=>x"00060",
2863=>x"00060",
2864=>x"00060",
2865=>x"00060",
2866=>x"00060",
2867=>x"00060",
2868=>x"00060",
2869=>x"00060",
2870=>x"00060",
2871=>x"00060",
2872=>x"00060",
2873=>x"00060",
2874=>x"00060",
2875=>x"00060",
2876=>x"00060",
2877=>x"00060",
2878=>x"00060",
2879=>x"00060",
2880=>x"00060",
2881=>x"00060",
2882=>x"00060",
2883=>x"00060",
2884=>x"00060",
2885=>x"00060",
2886=>x"00060",
2887=>x"00060",
2888=>x"00060",
2889=>x"00060",
2890=>x"00060",
2891=>x"00060",
2892=>x"00060",
2893=>x"00060",
2894=>x"00060",
2895=>x"00060",
2896=>x"00060",
2897=>x"00060",
2898=>x"00060",
2899=>x"00060",
2900=>x"00060",
2901=>x"00060",
2902=>x"00060",
2903=>x"00060",
2904=>x"00060",
2905=>x"00060",
2906=>x"00060",
2907=>x"00060",
2908=>x"00060",
2909=>x"00060",
2910=>x"00060",
2911=>x"00060",
2912=>x"00060",
2913=>x"00060",
2914=>x"00060",
2915=>x"00060",
2916=>x"00060",
2917=>x"00060",
2918=>x"00060",
2919=>x"00060",
2920=>x"00060",
2921=>x"00060",
2922=>x"00060",
2923=>x"00060",
2924=>x"00060",
2925=>x"00060",
2926=>x"00060",
2927=>x"00060",
2928=>x"00060",
2929=>x"00060",
2930=>x"00060",
2931=>x"00060",
2932=>x"00060",
2933=>x"00060",
2934=>x"00060",
2935=>x"00060",
2936=>x"00060",
2937=>x"00060",
2938=>x"00060",
2939=>x"00060",
2940=>x"00060",
2941=>x"00060",
2942=>x"00060",
2943=>x"00060",
2944=>x"00060",
2945=>x"00060",
2946=>x"00060",
2947=>x"00060",
2948=>x"00060",
2949=>x"00060",
2950=>x"00060",
2951=>x"00060",
2952=>x"00060",
2953=>x"00060",
2954=>x"00060",
2955=>x"00060",
2956=>x"00060",
2957=>x"00060",
2958=>x"00060",
2959=>x"00060",
2960=>x"00060",
2961=>x"00060",
2962=>x"00060",
2963=>x"00060",
2964=>x"00060",
2965=>x"00060",
2966=>x"00060",
2967=>x"00060",
2968=>x"00060",
2969=>x"00060",
2970=>x"00060",
2971=>x"00060",
2972=>x"00060",
2973=>x"00060",
2974=>x"00060",
2975=>x"00060",
2976=>x"00060",
2977=>x"00060",
2978=>x"00060",
2979=>x"00060",
2980=>x"00060",
2981=>x"00060",
2982=>x"00060",
2983=>x"00060",
2984=>x"00060",
2985=>x"00060",
2986=>x"00060",
2987=>x"00060",
2988=>x"00060",
2989=>x"00060",
2990=>x"00060",
2991=>x"00060",
2992=>x"00060",
2993=>x"00060",
2994=>x"00060",
2995=>x"00060",
2996=>x"00060",
2997=>x"00060",
2998=>x"00060",
2999=>x"00060",
3000=>x"00060",
3001=>x"00060",
3002=>x"00060",
3003=>x"00060",
3004=>x"00060",
3005=>x"00060",
3006=>x"00060",
3007=>x"00060",
3008=>x"00060",
3009=>x"00060",
3010=>x"00060",
3011=>x"00060",
3012=>x"00060",
3013=>x"00060",
3014=>x"00060",
3015=>x"00060",
3016=>x"00060",
3017=>x"00060",
3018=>x"00060",
3019=>x"00060",
3020=>x"00060",
3021=>x"00060",
3022=>x"00060",
3023=>x"00060",
3024=>x"00060",
3025=>x"00060",
3026=>x"00060",
3027=>x"00060",
3028=>x"00060",
3029=>x"00060",
3030=>x"00060",
3031=>x"00060",
3032=>x"00060",
3033=>x"00060",
3034=>x"00060",
3035=>x"00060",
3036=>x"00060",
3037=>x"00060",
3038=>x"00060",
3039=>x"00060",
3040=>x"00060",
3041=>x"00060",
3042=>x"00060",
3043=>x"00060",
3044=>x"00060",
3045=>x"00060",
3046=>x"00060",
3047=>x"00060",
3048=>x"00060",
3049=>x"00060",
3050=>x"00060",
3051=>x"00060",
3052=>x"00060",
3053=>x"00060",
3054=>x"00060",
3055=>x"00060",
3056=>x"00060",
3057=>x"00060",
3058=>x"00060",
3059=>x"00060",
3060=>x"00060",
3061=>x"00060",
3062=>x"00060",
3063=>x"00060",
3064=>x"00060",
3065=>x"00060",
3066=>x"00060",
3067=>x"00060",
3068=>x"00060",
3069=>x"00060",
3070=>x"00060",
3071=>x"00060",
3072=>x"00061",
3073=>x"00061",
3074=>x"00061",
3075=>x"00061",
3076=>x"00061",
3077=>x"00061",
3078=>x"00061",
3079=>x"00061",
3080=>x"00061",
3081=>x"00061",
3082=>x"00061",
3083=>x"00061",
3084=>x"00061",
3085=>x"00061",
3086=>x"00061",
3087=>x"00061",
3088=>x"00061",
3089=>x"00061",
3090=>x"00061",
3091=>x"00061",
3092=>x"00061",
3093=>x"00061",
3094=>x"00061",
3095=>x"00061",
3096=>x"00061",
3097=>x"00061",
3098=>x"00061",
3099=>x"00061",
3100=>x"00061",
3101=>x"00061",
3102=>x"00061",
3103=>x"00061",
3104=>x"00061",
3105=>x"00061",
3106=>x"00061",
3107=>x"00061",
3108=>x"00061",
3109=>x"00061",
3110=>x"00061",
3111=>x"00061",
3112=>x"00061",
3113=>x"00061",
3114=>x"00061",
3115=>x"00061",
3116=>x"00061",
3117=>x"00061",
3118=>x"00061",
3119=>x"00061",
3120=>x"00061",
3121=>x"00061",
3122=>x"00061",
3123=>x"00061",
3124=>x"00061",
3125=>x"00061",
3126=>x"00061",
3127=>x"00061",
3128=>x"00061",
3129=>x"00061",
3130=>x"00061",
3131=>x"00061",
3132=>x"00061",
3133=>x"00061",
3134=>x"00061",
3135=>x"00061",
3136=>x"00061",
3137=>x"00061",
3138=>x"00061",
3139=>x"00061",
3140=>x"00061",
3141=>x"00061",
3142=>x"00061",
3143=>x"00061",
3144=>x"00061",
3145=>x"00061",
3146=>x"00061",
3147=>x"00061",
3148=>x"00061",
3149=>x"00061",
3150=>x"00061",
3151=>x"00061",
3152=>x"00061",
3153=>x"00061",
3154=>x"00061",
3155=>x"00061",
3156=>x"00061",
3157=>x"00061",
3158=>x"00061",
3159=>x"00061",
3160=>x"00061",
3161=>x"00061",
3162=>x"00061",
3163=>x"00061",
3164=>x"00061",
3165=>x"00061",
3166=>x"00061",
3167=>x"00061",
3168=>x"00061",
3169=>x"00061",
3170=>x"00061",
3171=>x"00061",
3172=>x"00061",
3173=>x"00061",
3174=>x"00061",
3175=>x"00061",
3176=>x"00061",
3177=>x"00061",
3178=>x"00061",
3179=>x"00061",
3180=>x"00061",
3181=>x"00061",
3182=>x"00061",
3183=>x"00061",
3184=>x"00061",
3185=>x"00061",
3186=>x"00061",
3187=>x"00061",
3188=>x"00061",
3189=>x"00061",
3190=>x"00061",
3191=>x"00061",
3192=>x"00061",
3193=>x"00061",
3194=>x"00061",
3195=>x"00061",
3196=>x"00061",
3197=>x"00061",
3198=>x"00061",
3199=>x"00061",
3200=>x"00061",
3201=>x"00061",
3202=>x"00061",
3203=>x"00061",
3204=>x"00061",
3205=>x"00061",
3206=>x"00061",
3207=>x"00061",
3208=>x"00061",
3209=>x"00061",
3210=>x"00061",
3211=>x"00061",
3212=>x"00061",
3213=>x"00061",
3214=>x"00061",
3215=>x"00061",
3216=>x"00061",
3217=>x"00061",
3218=>x"00061",
3219=>x"00061",
3220=>x"00061",
3221=>x"00061",
3222=>x"00061",
3223=>x"00061",
3224=>x"00061",
3225=>x"00061",
3226=>x"00061",
3227=>x"00061",
3228=>x"00061",
3229=>x"00061",
3230=>x"00061",
3231=>x"00061",
3232=>x"00061",
3233=>x"00061",
3234=>x"00061",
3235=>x"00061",
3236=>x"00061",
3237=>x"00061",
3238=>x"00061",
3239=>x"00061",
3240=>x"00061",
3241=>x"00061",
3242=>x"00061",
3243=>x"00061",
3244=>x"00061",
3245=>x"00061",
3246=>x"00061",
3247=>x"00061",
3248=>x"00061",
3249=>x"00061",
3250=>x"00061",
3251=>x"00061",
3252=>x"00061",
3253=>x"00061",
3254=>x"00061",
3255=>x"00061",
3256=>x"00061",
3257=>x"00061",
3258=>x"00061",
3259=>x"00061",
3260=>x"00061",
3261=>x"00061",
3262=>x"00061",
3263=>x"00061",
3264=>x"00061",
3265=>x"00061",
3266=>x"00061",
3267=>x"00061",
3268=>x"00061",
3269=>x"00061",
3270=>x"00061",
3271=>x"00061",
3272=>x"00061",
3273=>x"00061",
3274=>x"00061",
3275=>x"00061",
3276=>x"00061",
3277=>x"00061",
3278=>x"00061",
3279=>x"00061",
3280=>x"00061",
3281=>x"00061",
3282=>x"00061",
3283=>x"00061",
3284=>x"00061",
3285=>x"00061",
3286=>x"00061",
3287=>x"00061",
3288=>x"00061",
3289=>x"00061",
3290=>x"00061",
3291=>x"00061",
3292=>x"00061",
3293=>x"00061",
3294=>x"00061",
3295=>x"00061",
3296=>x"00061",
3297=>x"00061",
3298=>x"00061",
3299=>x"00061",
3300=>x"00061",
3301=>x"00061",
3302=>x"00061",
3303=>x"00061",
3304=>x"00061",
3305=>x"00061",
3306=>x"00061",
3307=>x"00061",
3308=>x"00061",
3309=>x"00061",
3310=>x"00061",
3311=>x"00061",
3312=>x"00061",
3313=>x"00061",
3314=>x"00061",
3315=>x"00061",
3316=>x"00061",
3317=>x"00061",
3318=>x"00061",
3319=>x"00061",
3320=>x"00061",
3321=>x"00061",
3322=>x"00061",
3323=>x"00061",
3324=>x"00061",
3325=>x"00061",
3326=>x"00061",
3327=>x"00061",
3328=>x"00061",
3329=>x"00061",
3330=>x"00061",
3331=>x"00061",
3332=>x"00061",
3333=>x"00061",
3334=>x"00061",
3335=>x"00061",
3336=>x"00061",
3337=>x"00061",
3338=>x"00061",
3339=>x"00061",
3340=>x"00061",
3341=>x"00061",
3342=>x"00061",
3343=>x"00061",
3344=>x"00061",
3345=>x"00061",
3346=>x"00061",
3347=>x"00061",
3348=>x"00061",
3349=>x"00061",
3350=>x"00061",
3351=>x"00061",
3352=>x"00061",
3353=>x"00061",
3354=>x"00061",
3355=>x"00061",
3356=>x"00061",
3357=>x"00061",
3358=>x"00061",
3359=>x"00061",
3360=>x"00061",
3361=>x"00061",
3362=>x"00061",
3363=>x"00061",
3364=>x"00061",
3365=>x"00061",
3366=>x"00061",
3367=>x"00061",
3368=>x"00061",
3369=>x"00061",
3370=>x"00061",
3371=>x"00061",
3372=>x"00061",
3373=>x"00061",
3374=>x"00061",
3375=>x"00061",
3376=>x"00061",
3377=>x"00061",
3378=>x"00061",
3379=>x"00061",
3380=>x"00061",
3381=>x"00061",
3382=>x"00061",
3383=>x"00061",
3384=>x"00061",
3385=>x"00061",
3386=>x"00061",
3387=>x"00061",
3388=>x"00061",
3389=>x"00061",
3390=>x"00061",
3391=>x"00061",
3392=>x"00061",
3393=>x"00061",
3394=>x"00061",
3395=>x"00061",
3396=>x"00061",
3397=>x"00061",
3398=>x"00061",
3399=>x"00061",
3400=>x"00061",
3401=>x"00061",
3402=>x"00061",
3403=>x"00061",
3404=>x"00061",
3405=>x"00061",
3406=>x"00061",
3407=>x"00061",
3408=>x"00061",
3409=>x"00061",
3410=>x"00061",
3411=>x"00061",
3412=>x"00061",
3413=>x"00061",
3414=>x"00061",
3415=>x"00061",
3416=>x"00061",
3417=>x"00061",
3418=>x"00061",
3419=>x"00061",
3420=>x"00061",
3421=>x"00061",
3422=>x"00061",
3423=>x"00061",
3424=>x"00061",
3425=>x"00061",
3426=>x"00061",
3427=>x"00061",
3428=>x"00061",
3429=>x"00061",
3430=>x"00061",
3431=>x"00061",
3432=>x"00061",
3433=>x"00061",
3434=>x"00061",
3435=>x"00061",
3436=>x"00061",
3437=>x"00061",
3438=>x"00061",
3439=>x"00061",
3440=>x"00061",
3441=>x"00061",
3442=>x"00061",
3443=>x"00061",
3444=>x"00061",
3445=>x"00061",
3446=>x"00061",
3447=>x"00061",
3448=>x"00061",
3449=>x"00061",
3450=>x"00061",
3451=>x"00061",
3452=>x"00061",
3453=>x"00061",
3454=>x"00061",
3455=>x"00061",
3456=>x"00061",
3457=>x"00061",
3458=>x"00061",
3459=>x"00061",
3460=>x"00061",
3461=>x"00061",
3462=>x"00061",
3463=>x"00061",
3464=>x"00061",
3465=>x"00061",
3466=>x"00061",
3467=>x"00061",
3468=>x"00061",
3469=>x"00061",
3470=>x"00061",
3471=>x"00061",
3472=>x"00061",
3473=>x"00061",
3474=>x"00061",
3475=>x"00061",
3476=>x"00061",
3477=>x"00061",
3478=>x"00061",
3479=>x"00061",
3480=>x"00061",
3481=>x"00061",
3482=>x"00061",
3483=>x"00061",
3484=>x"00061",
3485=>x"00061",
3486=>x"00061",
3487=>x"00061",
3488=>x"00061",
3489=>x"00061",
3490=>x"00061",
3491=>x"00061",
3492=>x"00061",
3493=>x"00061",
3494=>x"00061",
3495=>x"00061",
3496=>x"00061",
3497=>x"00061",
3498=>x"00061",
3499=>x"00061",
3500=>x"00061",
3501=>x"00061",
3502=>x"00061",
3503=>x"00061",
3504=>x"00061",
3505=>x"00061",
3506=>x"00061",
3507=>x"00061",
3508=>x"00061",
3509=>x"00061",
3510=>x"00061",
3511=>x"00061",
3512=>x"00061",
3513=>x"00061",
3514=>x"00061",
3515=>x"00061",
3516=>x"00061",
3517=>x"00061",
3518=>x"00061",
3519=>x"00061",
3520=>x"00061",
3521=>x"00061",
3522=>x"00061",
3523=>x"00061",
3524=>x"00061",
3525=>x"00061",
3526=>x"00061",
3527=>x"00061",
3528=>x"00061",
3529=>x"00061",
3530=>x"00061",
3531=>x"00061",
3532=>x"00061",
3533=>x"00061",
3534=>x"00061",
3535=>x"00061",
3536=>x"00061",
3537=>x"00061",
3538=>x"00061",
3539=>x"00061",
3540=>x"00061",
3541=>x"00061",
3542=>x"00061",
3543=>x"00061",
3544=>x"00061",
3545=>x"00061",
3546=>x"00061",
3547=>x"00061",
3548=>x"00061",
3549=>x"00061",
3550=>x"00061",
3551=>x"00061",
3552=>x"00061",
3553=>x"00061",
3554=>x"00061",
3555=>x"00061",
3556=>x"00061",
3557=>x"00061",
3558=>x"00061",
3559=>x"00061",
3560=>x"00061",
3561=>x"00061",
3562=>x"00061",
3563=>x"00061",
3564=>x"00061",
3565=>x"00061",
3566=>x"00061",
3567=>x"00061",
3568=>x"00061",
3569=>x"00061",
3570=>x"00061",
3571=>x"00061",
3572=>x"00061",
3573=>x"00061",
3574=>x"00061",
3575=>x"00061",
3576=>x"00061",
3577=>x"00061",
3578=>x"00061",
3579=>x"00061",
3580=>x"00061",
3581=>x"00061",
3582=>x"00061",
3583=>x"00061",
3584=>x"00061",
3585=>x"00061",
3586=>x"00061",
3587=>x"00061",
3588=>x"00061",
3589=>x"00061",
3590=>x"00061",
3591=>x"00061",
3592=>x"00061",
3593=>x"00061",
3594=>x"00061",
3595=>x"00061",
3596=>x"00061",
3597=>x"00061",
3598=>x"00061",
3599=>x"00061",
3600=>x"00061",
3601=>x"00061",
3602=>x"00061",
3603=>x"00061",
3604=>x"00061",
3605=>x"00061",
3606=>x"00061",
3607=>x"00061",
3608=>x"00061",
3609=>x"00061",
3610=>x"00061",
3611=>x"00061",
3612=>x"00061",
3613=>x"00061",
3614=>x"00061",
3615=>x"00061",
3616=>x"00061",
3617=>x"00061",
3618=>x"00061",
3619=>x"00061",
3620=>x"00061",
3621=>x"00061",
3622=>x"00061",
3623=>x"00061",
3624=>x"00061",
3625=>x"00061",
3626=>x"00061",
3627=>x"00061",
3628=>x"00061",
3629=>x"00061",
3630=>x"00061",
3631=>x"00061",
3632=>x"00061",
3633=>x"00061",
3634=>x"00061",
3635=>x"00061",
3636=>x"00061",
3637=>x"00061",
3638=>x"00061",
3639=>x"00061",
3640=>x"00061",
3641=>x"00061",
3642=>x"00061",
3643=>x"00061",
3644=>x"00061",
3645=>x"00061",
3646=>x"00061",
3647=>x"00061",
3648=>x"00061",
3649=>x"00061",
3650=>x"00061",
3651=>x"00061",
3652=>x"00061",
3653=>x"00061",
3654=>x"00061",
3655=>x"00061",
3656=>x"00061",
3657=>x"00061",
3658=>x"00061",
3659=>x"00061",
3660=>x"00061",
3661=>x"00061",
3662=>x"00061",
3663=>x"00061",
3664=>x"00061",
3665=>x"00061",
3666=>x"00061",
3667=>x"00061",
3668=>x"00061",
3669=>x"00061",
3670=>x"00061",
3671=>x"00061",
3672=>x"00061",
3673=>x"00061",
3674=>x"00061",
3675=>x"00061",
3676=>x"00061",
3677=>x"00061",
3678=>x"00061",
3679=>x"00061",
3680=>x"00061",
3681=>x"00061",
3682=>x"00061",
3683=>x"00061",
3684=>x"00061",
3685=>x"00061",
3686=>x"00061",
3687=>x"00061",
3688=>x"00061",
3689=>x"00061",
3690=>x"00061",
3691=>x"00061",
3692=>x"00061",
3693=>x"00061",
3694=>x"00061",
3695=>x"00061",
3696=>x"00061",
3697=>x"00061",
3698=>x"00061",
3699=>x"00061",
3700=>x"00061",
3701=>x"00061",
3702=>x"00061",
3703=>x"00061",
3704=>x"00061",
3705=>x"00061",
3706=>x"00061",
3707=>x"00061",
3708=>x"00061",
3709=>x"00061",
3710=>x"00061",
3711=>x"00061",
3712=>x"00061",
3713=>x"00061",
3714=>x"00061",
3715=>x"00061",
3716=>x"00061",
3717=>x"00061",
3718=>x"00061",
3719=>x"00061",
3720=>x"00061",
3721=>x"00061",
3722=>x"00061",
3723=>x"00061",
3724=>x"00061",
3725=>x"00061",
3726=>x"00061",
3727=>x"00061",
3728=>x"00061",
3729=>x"00061",
3730=>x"00061",
3731=>x"00061",
3732=>x"00061",
3733=>x"00061",
3734=>x"00061",
3735=>x"00061",
3736=>x"00061",
3737=>x"00061",
3738=>x"00061",
3739=>x"00061",
3740=>x"00061",
3741=>x"00061",
3742=>x"00061",
3743=>x"00061",
3744=>x"00061",
3745=>x"00061",
3746=>x"00061",
3747=>x"00061",
3748=>x"00061",
3749=>x"00061",
3750=>x"00061",
3751=>x"00061",
3752=>x"00061",
3753=>x"00061",
3754=>x"00061",
3755=>x"00061",
3756=>x"00061",
3757=>x"00061",
3758=>x"00061",
3759=>x"00061",
3760=>x"00061",
3761=>x"00061",
3762=>x"00061",
3763=>x"00061",
3764=>x"00061",
3765=>x"00061",
3766=>x"00061",
3767=>x"00061",
3768=>x"00061",
3769=>x"00061",
3770=>x"00061",
3771=>x"00061",
3772=>x"00061",
3773=>x"00061",
3774=>x"00061",
3775=>x"00061",
3776=>x"00061",
3777=>x"00061",
3778=>x"00061",
3779=>x"00061",
3780=>x"00061",
3781=>x"00061",
3782=>x"00061",
3783=>x"00061",
3784=>x"00061",
3785=>x"00061",
3786=>x"00061",
3787=>x"00061",
3788=>x"00061",
3789=>x"00061",
3790=>x"00061",
3791=>x"00061",
3792=>x"00061",
3793=>x"00061",
3794=>x"00061",
3795=>x"00061",
3796=>x"00061",
3797=>x"00061",
3798=>x"00061",
3799=>x"00061",
3800=>x"00061",
3801=>x"00061",
3802=>x"00061",
3803=>x"00061",
3804=>x"00061",
3805=>x"00061",
3806=>x"00061",
3807=>x"00061",
3808=>x"00061",
3809=>x"00061",
3810=>x"00061",
3811=>x"00061",
3812=>x"00061",
3813=>x"00061",
3814=>x"00061",
3815=>x"00061",
3816=>x"00061",
3817=>x"00061",
3818=>x"00061",
3819=>x"00061",
3820=>x"00061",
3821=>x"00061",
3822=>x"00061",
3823=>x"00061",
3824=>x"00061",
3825=>x"00061",
3826=>x"00061",
3827=>x"00061",
3828=>x"00061",
3829=>x"00061",
3830=>x"00061",
3831=>x"00061",
3832=>x"00061",
3833=>x"00061",
3834=>x"00061",
3835=>x"00061",
3836=>x"00061",
3837=>x"00061",
3838=>x"00061",
3839=>x"00061",
3840=>x"00061",
3841=>x"00061",
3842=>x"00061",
3843=>x"00061",
3844=>x"00061",
3845=>x"00061",
3846=>x"00061",
3847=>x"00061",
3848=>x"00061",
3849=>x"00061",
3850=>x"00061",
3851=>x"00061",
3852=>x"00061",
3853=>x"00061",
3854=>x"00061",
3855=>x"00061",
3856=>x"00061",
3857=>x"00061",
3858=>x"00061",
3859=>x"00061",
3860=>x"00061",
3861=>x"00061",
3862=>x"00061",
3863=>x"00061",
3864=>x"00061",
3865=>x"00061",
3866=>x"00061",
3867=>x"00061",
3868=>x"00061",
3869=>x"00061",
3870=>x"00061",
3871=>x"00061",
3872=>x"00061",
3873=>x"00061",
3874=>x"00061",
3875=>x"00061",
3876=>x"00061",
3877=>x"00061",
3878=>x"00061",
3879=>x"00061",
3880=>x"00061",
3881=>x"00061",
3882=>x"00061",
3883=>x"00061",
3884=>x"00061",
3885=>x"00061",
3886=>x"00061",
3887=>x"00061",
3888=>x"00061",
3889=>x"00061",
3890=>x"00061",
3891=>x"00061",
3892=>x"00061",
3893=>x"00061",
3894=>x"00061",
3895=>x"00061",
3896=>x"00061",
3897=>x"00061",
3898=>x"00061",
3899=>x"00061",
3900=>x"00061",
3901=>x"00061",
3902=>x"00061",
3903=>x"00061",
3904=>x"00061",
3905=>x"00061",
3906=>x"00061",
3907=>x"00061",
3908=>x"00061",
3909=>x"00061",
3910=>x"00061",
3911=>x"00061",
3912=>x"00061",
3913=>x"00061",
3914=>x"00061",
3915=>x"00061",
3916=>x"00061",
3917=>x"00061",
3918=>x"00061",
3919=>x"00061",
3920=>x"00061",
3921=>x"00061",
3922=>x"00061",
3923=>x"00061",
3924=>x"00061",
3925=>x"00061",
3926=>x"00061",
3927=>x"00061",
3928=>x"00061",
3929=>x"00061",
3930=>x"00061",
3931=>x"00061",
3932=>x"00061",
3933=>x"00061",
3934=>x"00061",
3935=>x"00061",
3936=>x"00061",
3937=>x"00061",
3938=>x"00061",
3939=>x"00061",
3940=>x"00061",
3941=>x"00061",
3942=>x"00061",
3943=>x"00061",
3944=>x"00061",
3945=>x"00061",
3946=>x"00061",
3947=>x"00061",
3948=>x"00061",
3949=>x"00061",
3950=>x"00061",
3951=>x"00061",
3952=>x"00061",
3953=>x"00061",
3954=>x"00061",
3955=>x"00061",
3956=>x"00061",
3957=>x"00061",
3958=>x"00061",
3959=>x"00061",
3960=>x"00061",
3961=>x"00061",
3962=>x"00061",
3963=>x"00061",
3964=>x"00061",
3965=>x"00061",
3966=>x"00061",
3967=>x"00061",
3968=>x"00061",
3969=>x"00061",
3970=>x"00061",
3971=>x"00061",
3972=>x"00061",
3973=>x"00061",
3974=>x"00061",
3975=>x"00061",
3976=>x"00061",
3977=>x"00061",
3978=>x"00061",
3979=>x"00061",
3980=>x"00061",
3981=>x"00061",
3982=>x"00061",
3983=>x"00061",
3984=>x"00061",
3985=>x"00061",
3986=>x"00061",
3987=>x"00061",
3988=>x"00061",
3989=>x"00061",
3990=>x"00061",
3991=>x"00061",
3992=>x"00061",
3993=>x"00061",
3994=>x"00061",
3995=>x"00061",
3996=>x"00061",
3997=>x"00061",
3998=>x"00061",
3999=>x"00061",
4000=>x"00061",
4001=>x"00061",
4002=>x"00061",
4003=>x"00061",
4004=>x"00061",
4005=>x"00061",
4006=>x"00061",
4007=>x"00061",
4008=>x"00061",
4009=>x"00061",
4010=>x"00061",
4011=>x"00061",
4012=>x"00061",
4013=>x"00061",
4014=>x"00061",
4015=>x"00061",
4016=>x"00061",
4017=>x"00061",
4018=>x"00061",
4019=>x"00061",
4020=>x"00061",
4021=>x"00061",
4022=>x"00061",
4023=>x"00061",
4024=>x"00061",
4025=>x"00061",
4026=>x"00061",
4027=>x"00061",
4028=>x"00061",
4029=>x"00061",
4030=>x"00061",
4031=>x"00061",
4032=>x"00061",
4033=>x"00061",
4034=>x"00061",
4035=>x"00061",
4036=>x"00061",
4037=>x"00061",
4038=>x"00061",
4039=>x"00061",
4040=>x"00061",
4041=>x"00061",
4042=>x"00061",
4043=>x"00061",
4044=>x"00061",
4045=>x"00061",
4046=>x"00061",
4047=>x"00061",
4048=>x"00061",
4049=>x"00061",
4050=>x"00061",
4051=>x"00061",
4052=>x"00061",
4053=>x"00061",
4054=>x"00061",
4055=>x"00061",
4056=>x"00061",
4057=>x"00061",
4058=>x"00061",
4059=>x"00061",
4060=>x"00061",
4061=>x"00061",
4062=>x"00061",
4063=>x"00061",
4064=>x"00061",
4065=>x"00061",
4066=>x"00061",
4067=>x"00061",
4068=>x"00061",
4069=>x"00061",
4070=>x"00061",
4071=>x"00061",
4072=>x"00061",
4073=>x"00061",
4074=>x"00061",
4075=>x"00061",
4076=>x"00061",
4077=>x"00061",
4078=>x"00061",
4079=>x"00061",
4080=>x"00061",
4081=>x"00061",
4082=>x"00061",
4083=>x"00061",
4084=>x"00061",
4085=>x"00061",
4086=>x"00061",
4087=>x"00061",
4088=>x"00061",
4089=>x"00061",
4090=>x"00061",
4091=>x"00061",
4092=>x"00061",
4093=>x"00061",
4094=>x"00061",

others=>x"00000"
);
begin
Cout<=memory(to_integer(unsigned(addr)));

end Behavioral;